��   �E�A��*SYST�EM*��V9.3�0146 5/�27/2021 A   ����DCSS_C�PC_T  �4 $COMM�ENT $�ENABLE � $MODJG�RP_NUMKL�\  $U�FRM\] _VT�X M �   �$Y�Z1K �$Z2�STOP�_TYPKDSB�IO�IDXKE�NBL_CALM�D�USE_PR�EDIC? �EL�AY_TIMJS�PEED_CTR�LKOVR_LI�M? p D� L�0��UTOOi��O^ �x&S. � 8J\TC�u
!���0\� jY�0  � �C�HG_SIZ��$AP!�E�D�IS�]$!�C�_+{#s%O#J�p 	]$Jd#� �&s"�"{#p�)�$�'�_SE_EXPAN#N�{  ,$STAT/� DFP_B�ASE $�0K$4!� .6_�V7>H73
6J-� � }�\A�XS\UP�L�W�7��� �9`d4r �< w? �?�?��?�?�//�	7ELEM/ �T �&B.2NO0�G]@%CNHA�DF#~� $DATA)q
6e0  P�J�@ 2 
:&P5 �� 1�U*n   _VS iSZbRj0jR(�VyT�(�R%S{TROBOT�X�SARo�U~�V$CUR_���R4SETU4"	� $d P_�MGN�INP_ASSe#�PB!�  `CiH�77`e�.fXc�1�CONFIG�_CHK`E_PO|* }dSHRST�g�M^#/eOTHER7RBT�j_G]�R��dTv �ku�dVA�LD_7h�e�4HVT1r
0R HLHt� 0  lt<Ner�RFYhH~t�5�1ȕ ��W�_A$�Rd�TPH/ (G%Q�Q�Q�3?wBOX/ 8�@F!�F!�G �r���zTUIRi@ � ,�F�pE}R%@2 $�po l�_Sf��A�ZN/ 0 IF(@�p��Z_�0�_�0?wu0  @�QWyv	*���~ �$$CL�`  ����!���Q��Q�VE�RSION��  1b��$' 2 ?�Q  (�r����&@"�o��P���������������Ԓd��Cz   2����C���n����� ����ȟݯ���"� 4�F�H�j������֯ ǿ�������0�B� T�f�hύϜ�����ҿ ���ϐ��,�>�P�� tωߘϪ�d������� ��(�:�`�^�p߅� �߸��������� $�6�H�Z�o�~���� ��������� �2� D�j�Xz�������� ����.@R dy������ �	//*<N�b/ ��/����/�? ?&/8/J/\/n/�?�/ �?�/�/�?�/OO%O 4?F?X?j?lO�?�O�? �?�?�O�O_!_0OBO TOfOxO�O�_�_�O�O �_�Ooo�_>_P_b_ t_/o�_�o�_�_�o�_ �o+:oLo^o�o�o �o�4�o�o� � '�6HZl~��� ���������#�5� D�V�h���|����� ԏ���
��1�@�R� d�v���������П� ����-�?�N�`�r� �������̯ޯ�� �)�;�J�\�n����� �϶���ڿ���%� 7�I�X�j�|ώϐ߲� ����������3�E� T�f�xߊߜ߮߰��� ������/�A���b� t���S��������� ���=O^�p��� �������X��  $9KZl~�� ������ !/ G/Y/hz���/� �/��
/?./C?U? d/v/�/�/�/�?�/�? �/?O*??OQOcOr? �?�?<O�O�?�O�?O O)_8OM___nO�O�O �O�O�_�O�_�O_%o 4_Io[omo|_�_�_�_ �o�_�o�_oBo3" Wixo�o�o�o�o�o ��/�>S�e� �����w���� ��Џ:�,�a�s��������̏ʏ܋�$D�CSS_CSC �2���?Q  P����<�މd�m�0��� T���x�ٯ����ү 3���W��{�>���b� ��տ��������A� �e�w�:ϛ�^Ͽς� �Ϧ������=� �a� $߅�Hߩ�l߹��ߢ� ���'���K��o�2� ���h�������GRP 2�� ����	ԟU�@� y�d������������� 	��?*cN� r������ M8q\�� ����/�/7/ "/[/F//j/�/�/�/ �/�/�/?�/?E?0? i?T?�?�?�?|?�?�? �?�?	O/OOSO>OwO �O�OfO�O�O�O�O_ �O_=_(_a_s_�_P_ �_�_�_�_�_�_o'o�oKo�_GSTA�T 2��'���< ��5-�A?1Ԍ>���>ER	<k��_?{,�?.�?8˾~�_D�(�Ĳ��1DYh��:`<��e?}������3;��4���?�  �a���`4��ZC�y�Ĺ�����f�Z��=�Nn?�{п 8=�j7�\���i��U�ĩ���D�y=�q����X�?~�X>©�`�����(�{�>���=��;���ĪC]D�?�$y>_�?|���Q�bpfp�jp>��=�2�?}�JD�ĸ�ȿ/�D
��z8��?0�=>�������2��}I�.w��`>~� �o�o�o�b�f�`މ:��Ĵ�&�m��z� ����n���ʏ���jK� ��0h.��6��>�l� R�d����������П � ���:�h����� �������֏�r�� J�$�R�8�J���n��� ��п��ؿ����<� "�4�Vτφ����ϼ������p�����6�:���*��;�>��Ͻ�F[��� =�F����A�7ώ���C� "Y�m<;�C���7a4����1wx��arѼ�o��a@e������m�"�?�]ߍ>�[]���}�>�W��]�J����q��'1D	��y;�X�R��D?z��?s�<�;�����I��7��?z}k>�R����{��2�,D=�����W�R�?z�ɼ7�s�����MY��;�F/AM}���y�C���y<I)��߾�F�.�<�MY���C�;�� �F��? O�G�)�;�M�oϑ�S��x���"��� X�j������Ϭ��� ��������H. `~dv���� ��L�>P*t� |������  /.//6/d/J/\/~/ �/�/�/�/�/�/?�/ hZ?l?F?�?�?|?�� ��R�d�v߈ߚ߬߾� ��������*�<�N� `�r��O�?�?�??.? ��B?�?�_�?�_�_o ��_0o>?HofoLo^o �o�o�o�o�o�o�o  4bHj�~ �_����"�o� L��D�f���z���ʏ ��ҏ �����H�.� P�~�d���������� ��,�>��6_H_�?  OO$O6OHOZOlO~O �O�O�O�O�O�O�O_ ��b�t�����ʟ�_ޟ L�Z�P�FϐϢ�<�"� ��ڟ��������J� 0�R߀�fߘ߶ߜ߮� �������4���v� ��b����>���R� ���0��8�f�L�n� ��������������  "P6���~ ���ҿ俊����� ��ү�����,�>� P�b�t�������/� "Df(�z��/ ��/,?>?��/h?v �?�?�?�?�?�?�?�? OO4ORO8OJOlO�O �O�O�O�O ?_$_�O H_Z_P?�O�_�O|_�_ �_�_�_o�_
o8oo 0oRo�ofo�o�o�o�o �o�o<_.@dv Pn/�/&8J\n �������� /"/4/F/����� �o�/����~� ȟڟt_Z���:�  �2�T���h������� Я�ԯ��6��>� l�R������������ �v� ϊ��:�h�N� pϞτϦ��Ϻ����� ��$�R�8�Z߈�n� ؿ���߶� ����
� �����
��.� @�R�d�v��������� Џ�T�6�H�Z�|ߞ� `��� �.$�dv �����߸��� �&T:l� p�����/� XJ/\/6/�/�/�/ �/&/�/�/?�/?:?  ?B?p?V?h?�?�?�? �?�?�?�?$O
Ot/fO xORO�O�O�O����^� p�����������  ��$�6�H�Z�l�~� �_�O�O�OO:O��NO �O�o�O�o �/�o <JOTrXj�� �����&��� @�n�T�v������o� ��ҏ�.�$��X� P�r�������֟��ޟ ���&�T�:�\��� p������������8�J�X��$DCS�S_JPC 2�B�Q (G DOP������ ���`��ݿ������ ���[�*�i�Nϣ�r� �ϖ��Ϻ����3�� �i�8�J�\߱߀��� ���������A��"� w�F�X�j������ ���+���O��0�r� ��f�x��������� ��9],�P� t�����#� 1k:�^�� �����1/ // $/y/H/�/l/�/�/�/ �/	?�/�/??? ?2? �?V?�?z?�?�?�?�? O�?�?:O_O.O@O�O dOvO�O�O�O_�O%_ �OI__m_<_N_�_r_��_�_�_�_�_�cj�S
s�w�L�_Woo{o�`dFo�ojo�o�o�o �o�o3�oW{ BTf����� ��A��e�,���P� ��t���������Ώ�� �O��s�:���^��� ��ߟ���ʟ'�� � �[���H���l�ɯ�� ���د5���Y� � g�D���h�z������� ¿��C�
�g�.ϋ� Rϯ�v��ϚϬϾ�� -���Q��u�<ߙ�`� �߄��ߨ������� M��&�8�J��n��� ��������7���[� "��F�X�j������� ����!��Ei0 �T�x���� ���Sw>� b����/�(d�MODEL 2�5kx��
 �<�c(  �|(�/i/{/�/ �/�/�/�/�/�/F?? /?|?S?e?w?�?�?�? �?�?�?0OOO+O=O OOaO�_�O[/�O�O_ �O�O>__'_9_�_]_ o_�_�_�_�_�_�_�_ :oo#opoGoYo�o}o �o�o�o�o�o�O�O�O �o~�ogy�� ����2�	��-� ?�Q�c�������揽� Ϗ����d�;�M� ��5Gu�����o�ݟ ���%�r�I�[��� �������ǯٯ&��� �\�3�E�W�i�{��� ڿ��ÿϫ������ j��S�eϲωϛ��� ���������f�=� Oߜ�s߅��ߩ߻��� ����P�'�9��!� 3�E�s��[�����(� ���^�5�G�Y�k�}� ������������ 1C�gy�� ���� ����� ?Q�u���� ���/R/)/;/�/ _/q/�/�/�/�/?�/ �/<??%?7?�?1 _?q?�?�?�?O�?�? JO!O3OEO�OiO{O�O �O�O�O�O�O�OF__ /_|_S_e_�_�_�_�_ �?o�?�_�_To+o=o �oaoso�o�o�o�o �o�o>'9K] o������� ��#��_��oK�]� ʏ���� �׏���� �1�~�U�g������� ����ӟ�2�	��h� ?�Q�c�u�����o��� ����ӯ@��)�v�M� _�q���������˿ݿ *���%�r�I�[Ϩ� ϑ��ϵ�����&��� ����	�7�I߶�1� �߱�������4��� j�A�S�e�w����� ���������+�=� O���s�����m�߭� ��,��'9K] �������� �^5G�k} ����/��H/ ����#/5/�//�/�/ �/�/�/ ?�/	?V?-? ??Q?�?u?�?�?�?�? 
O�?�?ORO)O;O�O _OqO�OY/k/}/�O�O �O__`_7_I_�_m_ _�_�_�_�_o�_�_ Jo!o3oEoWoio{o�o �o�o�o�o�o�o�OX �O!3	w��� ������+�=� ��a�s���������͏ ߏ�>��'�t�K�]��o����$DCSS�_PSTAT ����Ց�Q    l��� � (��-��Q���v�  t�֐�������������Օ⯐�ׯ	�Ɣ�SETUP 	NՙBȘ����� :�T�Ϭu�d����������I�ƔT1SC �2
-�����Cz�����)��CP [R�D�DN tφ�@�ϼ��ϝ��� ����:�L�^�-߂� ��cߥ����߫� �� $���H�Z�l�;��� ��������� �2� �V�h�z�I������� ��������	.@ dv���`ϵ�N ���3EW& {��n���� //�A/S/e/4/�/ �/�/|/�/�/�/�/? +?�/?a?s?B?�?�? �?�?�?�?O�?'O9O KOOoO�OPO�O�O�O ��O�O_�O5_G_Y_ (_}_�_�_p_�_�_�_ �_oo�_CoUogo6o �o�o�o~o�o�o�o�o -�oQcuD� �������)� ;�
��q���R����� ˏ������O7�I� [�������r�ǟٟ �����!��E�W�i� 8���������կ篶� ȯ�/���S�e�w�F� ������������ֿ +�=��a�sυ�Tϩ� ���Ϝ�������9� K�]�,��ߓ��t��� �ߪ����#���G�Y� k�:��������� ����1� �U�g�y� H��������������� ��-?cu�V ������ ;Mq��d߹ ��d//%/�I/ [/m/</�/�/r/�/�/ �/�/?!?3??W?i? {?J?�?�?�?�?�?�? �?O/OAOOeOwO�O XO�O�O�O�O�O_�O �O=_O__s_�_�_f_ �_�_�_�oo'o�_ Ko]ooo>o�o�oto�o �o�o�o#5Y k}L����� ���1�C��g�y� ��Z�����ӏ����	� ؏-�?�Q� �u����� h���ϟ៰���)� �_M�_��@�����v� ˯ݯﯾ��%�7�� [�m��N�������ٿ ���̿!�3�E��i� {ύ�\ϱ��ϒϤ��� ���/�A�S�"�w߉� ��j߿����߲������=�O�a�0��$D�CSS_TCPM�AP  ������Q W@ 8�8�8�8���8�8��8�8�	8�
8��8�8�8�8��9�  8�8��8�8�8�8�R8�8�8�8�8�U8�8�8�8�U 8�!8�"8�#8�U$8�%8�&8�'8�U(8�)8�*8�+8�U,8�-8�.8�/8�U08�18�28�38�U48�58�68�78�U88�98�:8�;8�U<8�=8�>8�?8��@�UIRO 2]������� ������ $6H Zl~�������7���7�� [m����� ��/!/3/E/W/i/ {/�/�/<�/�/�/ ??/?A?S?e?w?�? �?�?�?�?�?�?OO �/=O�/aOsO�O�O�O �O�O�O�O__'_9_ K_]_o_�_�_�_0O�_�{�UIZN 2.��	 �����
o o.o4�o\ono�oCo �o�o�o�o�o�o�o 4FX'|��c ������0�B� �f�x�G�������ҏ �������>�P�b� %�������y�Ο��� ���(�:�	�^�p��� E�W���ʯ��� ����_��UFRM R.�����8;�h� z�9����Կ��� 
����@�R�-�vψ� cϬϾϙ�������� *�<�S�`�r�ߖߨ� �����߹�����8� J�%�n��[����� ��������"�4�K�X� j�	�����{������� ����BT/x �e������ ,C�Pb�� s����//� :/L/'/p/�/]/�/�/ �/�/�/�/?$?;2? Z?l?G?�?�?}?�?�? �?�?O�?2ODOOhO zOUO�O�O�O�O�O�O 
__3?E?R_d__�_ �_u_�_�_�_�_o�_ *o<oo`oroMo�o�o �o�o�o�o�o&=_ J\�o��m�� ����"�4��E� j�|�W�������֏� Ï��5B�T��x� ��e�������џ��� �,�>��b�t�O��� ����ί௻����