��  
J��A��*SYST�EM*��V9.3�0146 5/�27/2021 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP�fBI�IZ@���ALRM_RwECO"  � wALM�"ENB����&ON�!� MD�G/ 0 $?DEBUG1A�"d�$3AO� ."��!_IF� �� 
$ENABL�@C#� P dC#U5K�!MA�B �"�
� OG�f 0�CURR_D1P $�Q3LIN@S1I4$�C$AUSOd�A�PPINFOEQ�/ �L A �?1�5/ H ��79EQUI�P 2�0NA�M� ��2_OV�R�$VERS�I� � PCOU�PLE,   �$�!PPV1CES0�!H �1�2> �1�	 � $S�OFT�T_ID�BTOTAL_EeQ� Q1]@NO`B�U SPI_IND�E]uEXBSCR�EEN_�4BSIG�0O%KW@�PK_FI0�	$THKY�GP�ANEhD � D_UMMY1d�D��!U4 Q���A�RG1R�
 � _$TIT1d  ��� 7Td7T� 7TP�7T55V65V75V8
5V95W05W>W�A7UPRWQ7UfW1pW1zW�1�W1�W2�R�!S�BN_CF�!�0$!J� ; 
2��1_CMNT�?$FLAGS]��CHE"$Nb_�OPT�2�� EL�LSETUP 7 `�0HO�0 �PRZ1%{cMAC{RO�bREPR�hD0D+t@��b{�e[HM MN�B
1^�0UTOB U��0 9DoEVIC4STI�0��� P@13��`B�Qdf"VAL�#IS�P_UNI�#p_�DOv7IyFR_F�@K%D13�;A�c�C_WA?t�a�z�OFF_@N�DEL�xLF0q�A�q�r?q�p�C?�`�A�E�C#�s�AsTB�t��MO� ��sE � [Mp�s��2�REV�gBILF�!XI� ~%�R  � �OD}`j�$kNO`M�Qb�x�/�"u�� ������!X�@Dd� p E RD_�Eb��$FSS�B�&W`KBD_S�E2uAG� G�2B "_��B�� V�t�:5`ׁQCe`�a_E�Du � � �C2��`S�p�4%y$l �t$OP�@rQB�qy�_OK���0, P_C� y��dxh�U �`LACI�!��a���� FqCOsMM� �0$D���ϑ�@�pX��OR BIGALLOW�G (KD2�2�@VAR5�d!�AB �`�BL[@S � ,�KJqM�H`S�pZ@M�_O]z���C�Fd X�0GR�@��M�NFL�I���;@UIRE�84�"� SWIT�=$/0_No`S�"C�F_�G� �>0WARNMxp�d��%`LI�V`NS]T� COR-r�FLTR�TRA�T T�`� $A�CCqS�� X�r�$ORI�.&ӧR�T�`_SFgPC�HGV0I�p�T���PA�I��T�撡HK�� �� �#@a���HD)R�B��2�BJ; �CT��3�4�5�U6�7�8�9>�x��x@�2 @� TRQ��$%f��ր����_U�����`{COc <� �����Ȩ3�2��LL�ECM�-�MUL�TIV4�"$��A
2FS�ILDD�
1��z@T_1b  4� STY2�b4�=@�)24����E��� |9$��.p���6�I`�* \�T�O��E��EXT����ї��B�ў22��0D��@`��1b.'�B �G�Q� �"Q�/%�ap��X�%�?sONLCՂU� Sҟ�;A�Ɨ�M8�� � CՋO�! L�0a�� �X׻pAβ$JOB`B�������IGO�" dӀ�����X��-'x���G�ҧ@�_M\��b# tӀF� f�CNG�AiBA�  ϑ��!���/1��À�0����R0P/p����$
�|��BqhF]�
2J]�_RN���C`J`�e�J
?�D/5C�	�ӧ�� �@{  AzO3л!7% \�0RO�6�� �IT�s� NOM_8pn#�c �Ѭ�TU�@P� )� ��&+P��� bӨP�	ݭ��RAx@�n �3�A���
$TYF3%#D3
T�ԢwpU�13�}�%mH,rzT1�E� ��ޣ�#ݤ�%ߢQl�YNT�"� DBG�DE�!'D�]�P�U���@t����"��AqX��"�uTAI2s�BUFۆ��?!�1(c ��P&V`PI84�'mP�'M�(M��)B �&F�'SIMsQS�@ZKEE3PAT�zЙ8"�\"�!_MC��)SЌ0��`JB���ľaDECg:� g5.�����* �U�CHNS�_EMPͲ$G���7�_��c;�1g_FP)�TC�6S���5�`%��4�} �V����W��JR�����SEGFRA�q�Oaa #PT_LsIN�KCPVF�� �C$+���ckBZ���PBzrN4	,` +�ԦE��A�0� �Ad0o`Ar�D���Id1�SIZh���	T�FT`�C�Z1Y�ARSm� �CP@'�Ic\1@cX��0<@L����0�VC3RCߥ�sCC���U@1@�X�1��2�Mpq@�U�1`�X�Q�UDݤأiCk�p��
DK`0݀f��RhEVRf �UFha_	EF�0N�f �Pd1�&h��5��jC}�+�VSCA�[��A�f�2��4-2)��p��SFV�P�#t1BP�K2�4��.��	�ׇMARG����a�F@@���1D8cQ���0LEW�-��R�P<��o�lI2RɄ/������ȯ��� 5ڡR� HANC��$LG5��a�� Ӑ��ـF��Ae����0R�r�3@�����@�@ ;�RA��@�A�Z�0��N`�O��F#CT���p�F��R��0P0b ADI�O �a���a���&�ӄ5�5����S[�g���'BMPUD(PY�1���AESCPjc�WꍠN  Sh�XYZ'WPR�c�����	/����0  E�PI8���41��n@_C�$ϑW��N}U0MMENU�2)�TIT]q<�b�1%ECA:"Z_#`S3 ��� �!S�[v�NO_HEADE���c~���l�0��$ x��4.��RE�� "��4�4 T!�b�5CIGRTR�0�W�XL�t2,dC�gRJ��O��� ERRLd��5X�&Q/�OR�B$C��������$RUN_�O7��P$SYS�2�4i�/���!qV��dA *�PXWO�A`�6e@$SK�o�":!DBT�pT+RL�7.��P�����[�INDU DJ$�p�_�`�!������PL�A_2WA���E��D!�!�%Rh��UMMYi9f�H�1� 琓DB���8���!PR�Q 
����9���9 Ц$�r�$ Q�L���:�����P�;,��%�PC�<����WENEC0TNr=���%��COR��>�H mO�@79$LC�:$�ê"�{�T�R@�AUBb�_D��� ROS �"SKS��Zr���� =�����PA��JVBE�TURN���SMR�(�U #�CRr�E�WMDB0GNA9LV �"$LA� ��*;$P,p<$P���=�!�P1C2��PDO^@,s�o�Y��Rs�GO_AW���MO��pB��_�CSSҐSTCY��?�����0����ID���2��2
��NK�ON�J��v`�I~� @ P �$L�RB�B֓P�I��PO�I_B�Y�r�-�TVR��HwNDG7�A H�`�1	�@ݦDSBLIAN�y���0�昰��LS<BZ�0� f��FB���FE}�@������5<CK �$DO�1�C"�MC�0��4+��R�HɀWU0��w�6ELE�Lr����\ �DӠ$�г�INQK$���U��L�cHA��Q{P$�#�{P���VE ��˰MDLy 2AD0����)C��J{R6 {R<YO�����0x����SLAVNrFxBINS ,��#,�X��`��GrC��\�   UL�����SHOWF!HF[3BT�!���&�&r��I�@,$\`�p���
�%
�,�u2�FI�g"���f#ID׀c&�c&W9RՓ�"NTVh"sVEԔ2�SKI3�lA�C;3�'2UB�1Jp�f�1��
DSAF���#7_SVl�EXC�LUձY��rON	L�0K3Y�Ȁ^�HI_V��RPPkLY�RysHIX �_&y3_M�b��VORFY_�w2M�s_$IOCt�OՓD�1�P1UB�43O�F|5LS��N�Q�47�I�2��:@ðP��i$���6A� CNr@�N�AE��&C���GCH	D�y�_����%0}�CP�#aDT)�x�NB_VAL:�9�H#���� JЪ�TqAа_��� ��J� CLtK��pT�ЂU� ^G�D��p���?L D $ۀx�g�*S!}P3V_<0>\H<S�2p�s@K��M��Ӵrx�$R� L �S}G�` N �0�CUR�����S��Q������Њ��X���VANNUN��JE�S���PLY�
�&�ia���j0f�BEF2�I.��O @�`F�R��	$TOT �	�Q�@)�Q�C
Cf�KaM��NI��P��bU��b�Ab!�dDAYH�L�OAD�FėbG�5��cEF(pXI��Q��<�P�O�`�QU��_�QOqR"PP��Q�&pu2sE��;s�e� Q� �w!q	�� �A\�q)qS 0)a{q�i{qO��v�DU ��u���CA} TZb|��� �n�IDLE_PW�T��wtW�o�V�V�_vp� V��DIA�G��U� 1$�@Z ՓTߒw&�p�� ,�)�wR��au�VS���SW�c�[�3��pD�!u� R�y!qOH7u�qPPLS�wIR�wB�� �rTC��v*`ǂx����x w@����u� T�� &p��*�RQDW&��MS��&�A{���<Q�uLIFE�2cAPX��Nc�-�l�a$a�-�C��cC��0P�x�N��Y7���FLAwCaOV��x�O�|�wSUPPOаIA��_ٔ�U��C_Xj���r��Z�W����o��k�jҳXZ�uY2_�C"��T����+�N�`)��aN ��^Pv�BI{CTL$V `��CACHSرǣ��UT3�N� UFFI�g ��F���bG�6�b�aMSWW 8`KEYoIMAG��TMW� �cE��RA����p �VIEm���X ��BGL�$`�#?G� 	��@��Y"PmE ST9�!�� I���7��� ���`��EMAI� �ѤA-�^~AFAUL��Z}��ӤB� ~�U� h��STB.`N#[3�R����к�h6�@�#��LD�EBU���~�T�2�)q\< $di�Svp�pIT3�BUFڧ�!ڧ��N�f1g�SUB���C��$��j¯���SAV �Ţ�'�~���w���_0rfP��ORDn��y�_���ũA=�OT(��V �sP�0M�%fԌ�Bc�AX�M`�0Xؕ�-3�_Gc�
A��DYN_���`]� <0pD�������M�r��T@F�p��g@DI�A��EDT_k�� �a^$�m0G��ha&�SU����k���� F~� 7_ ( SV|������!zi�2�T`� ��0�D�7C_Rx�IKp����R��R=����2�'DSPU�k�P��IM������E2�@�U��ΐW���M��I�P�#k㡁����TH�}����pT{���H9S�ӧ�BSC�$����pVy�s��{�_�D�CONV71G �{�}����Fc��ad���Њ�q�SC���}�MERr42�F�BCMPr31�ETnf a3�FU�DU��[AO0U�=B�CD��E�W�	��`O�`��b.s�Qs�q�Q� s��AMSwAQ
�@�T ����b ��ac�� "�pp���$ZO(��B���@U��JD�P�$�CN��C�@��GRO�U�� r�xSɠ�CMN�nnnr��H �S���CYC������a>1	*DEp1_D뢧pRO�T�v�`��0OaR&ncQ' 	$:�[�%�%�W��@&�!AL`��ad�Bi��A<Cj�p@B��Ph��R�@TV�ge ,@{P�!'զ!��i�L���1d 
�v�NOAA�af"R4�e4�e)P�A2C�@)5�#�b�2jо gH *)1L�0�n@q2 ��.`d@W�6�A�6A��6�a�6�a�6��67
�98�99�:c��8�:U1�:1�:1�:1�:U1�:1�:1�:1J�2J2�;�:2�:2��:2�:2�:2�:2��:2J3J3�:3T�;�:3�:3�:3�:U3�:3�:3J4B&]XT��ah��� ����������W�� ��FDR�iTu�VE�p_�f�#a,s�f�RE1F�1x��OVM��IeARiT7ROVRiDT��rjMX�lINRi��qjN	�IND�`Ir
�h��f���G��΃{`g �l�R�D6v{`RIVx ��x�GEAR��KIOI�KBbv�N��0xEFFRiC�a�>x�Z_MCMW�f�� �FϐURjx� (0��? ����?�pb�?�qE)��qg����b�k"��P}��R�I�0��ETUP?2_ l а��#TD3�)���Tb�qp�w�u��BAC��Gm T�����)��%) ~�"�qIFI�"v�M�00N��PT3�]FLUI�$�n � !P�k�URށѪ�� �s��Ne#EMP��$ʂ]S~�?xրJ�"�/�R�VRT�P�x/$SHOˁLH��ASS��]ђ�5��TBG_�3,��3,��3�,��3,��3FORC�
�`���o �F�Uyq1��|�2*�q���}�n�p |�`7NAV��ʀ����>`S���$VgISI�`�SCm�CSE�p�ZЉ2V& O�!$�'>`m �&�$� I#p����FMR2eq "bC��#a&� =�'g.@Rif�fe�Bb_1Q�nLIM�IT_Q�?C_L�M�f}DGCLF�c�aDY�Z��pB�d5�f�o�d�qM#��r`�� T��FS:С�s P��Pq�&�pp$EX_q���q�1�����jq�3��5���G���et ��`SW��ON�xc\�0�\��GeGRbp�U��B�KIO1l@ �`POy�*�� ���M�"Ox� SMz� E������`�� _E u x��a��TERMz�9v�� �ORI��}w��  �SM 	O�r�x��M�� ���y��m�UP^  �z� -�a�Quʀ���v��G��ELTO�� ����FI���yp��>�|���w$UFR;�$00�l�:��OTyת�TT#`��wNST�PATJ�=��PTHJ�8 �Eg J��8�ART�ѠA�8�Ѡ��D�REyL��I�SHFT<�(7ѧ���_�R 5J�� ��$��7�yС 7������ �I�ͤ�U�� A PAYLyO��DYN_����p��ќ�15G�ERV�0r���"��R������?Qj���1j�RC��q15ASYMFL3TR157�WJJ��Q��`E�s������;U�!������8�����P������Q�OR�ML:�� GRi�d{w���OƦ�f�� �9H�!v�| ԍ�n�,�:�OC0�4�$OP �����>a��RE���RN��с!�1��e��R��8��H�e$PWR�`#ݓ��R_����̐ D��UD�r����W� ]}�p$HG�!� �ADDR�Hl�G`������PRR��a~ H�PSSC �?S��3��3��3�SEe����HSC�D_MN�������%b!$ ��HO�L�!�R �U�V�C�RO��@ѯ�ND_�Ci2��v�GR'OUP����_�p��4���1�A,b��A� ?P�Ga��0��0���0,bA�!r��SAGVED�G#�T@�c� $� ��_!D�P7��AP� ��}t�HTTP_0�Ha� ('0OB�J�H�$�L�E���#v0� �� �W���P_�aT�_��"S��c㚈KR�Lj	HITCOU6a"��L�� �"�`Ɔ� l� SS�`��TJQUERY_�FLA��_WE�BSOC��HW�A=�a�� �IONCPU��̑O�6 1����0�1�1~iR �IOLN*��� 8�PR(�`�$SL��$INoPUT_H�$* bHP����0SLH 
a��0OLEHD���E��=IO{ F_�ASx��0�$LE��'E�'���|N�`��C��
Ct�HY�Wp�A�Ck�~AUOPu�� `�@�A��b�D�`�FQ< Pc�* 	W�-Q�F:R#Vt�IP_sME����� X�@cIP� ��lR_N���~0̱���S�V�Q�kSPH�� ]�!�B-G���ϐM�ᐁg� l��Z�TA��� A��TI3UM���y��U��PS�VBUy�IDi�$2��e `e��Rb���CB"�Zd�T@Nhhy��ie�IRCA_C}N�` � ��)mG@CY� EA�C �a呯lPc��gŃ�x�cW�DAY_$`hNTVA��3`wp;B��cwSCA��FwCL�$a��$b␐��Oopd��|e�uN_��Cp��`$b�a�P�CBn���q!Q�"�$`a �hn� 2�� �@�QH����p0��v�"�PLAB�Ѹ�y��UNI�����ITYS�Q�"URR���w������R_URL���$AUEN�3�̑� ��TT_UńA�BKY_T�\�!J4�0r��gP$���D灬0RUԀ��A��dFAށJb1�FL��䜀��
���
�U�JR��� �� F���P�΀e�)�DXsg$J7�ǒJ8T�!7Ȱ�b]�o�7�P�y8��S�APHI!��Q^���D��J7�J82�L_KE~A�  �K�0�LMra � <�opXR�@�0�cWA?TCH_VA���<[��&FIELzP�1y]pؒu�� ����1V|5�9�CTr�D�ڄU�pLD_��3 x·_M8��yDbq�LNTK��N]COOh ��N%�B��T1?�����JĦ�/��p��LGi���� $�iLG_SIZ�$��R�
�,�@
�FD�I	� � K��,�|�"��� �������@��7����|������/�_��_CM}�߱LP��AF����2(�B��,��,��@,�7�8�I+�B�[�`,�s�D�6��RS��6��  &�ZI���SN��LNH����@-&0DE�EMBǐ ��}��#����L����7DAU��EA� �0����GH����@�BOO���3 C�B`PITp3D��� �FRE�P[�SCR�3�AD@ �2�MARGINAm��@+F�C����-4�AS�#BW�ԓA�ĞCJG=M��MNCH��AFNΒ��K猀��UF$�y�$�FWDv$�HL[�STP$��V$�<�$�K�$�RS"��Hi�@�FC{�q�  �Ck ����U�!8�@�׌���N��C+�G��PO/�v��q����Q&�EX�GTUI�Ig��s�`g��" ���Ӯ��A�F"+ŐT w���w�N{�A�NA�BۤAVAIp���Qs��DCS�`P**O0O<�S��ZGSS��IGN �$p2��Z��qn3DEV��LL��#2�Dc�P�3�RaT.�$�I��2�dt�r�A�P �3��qp@�3i�PS1"2"3"��`�+ �P� ��+��٤EZ�Dek!n5J�XY�o��ST�@R��Y��� �$E�C�H�� ��8A@�P� L�0�O ���H�V�0�B�4� �B$0�u�_ �  �0�!=sx�p#�MB_PN��5��P�CC8�TRIqN���@BAS���ѩ&IRQ�&�1M�C��� �&�C�LDP�@��TRQ�LI:�Ȇ�)�$FL ���!�3OqD'�7Ƙ0LD5�$5OR�G΁��$2ԸRESERV�4p4�3p4�2<�$�� �s��$0���$5�PT� ��	T1�4�6RCLCMC�4p?�?�94�3��M���Ac�����MA}��`�sвU���T eEp�~Q�� F� i�� � ���HRS_RU���:!�tA�`��FgREQ�$��	�OVER
`2��Pt\.�P-�EFI+`#%!�t�
|C�4Ǣ \���Ao�$9Ub�r?s�$qPS!�	�C���4��R=S�3Us`HA?�(,@$L�MIS�C�� d��bR�Q�	�����`��V��XAX��Ӑ�W>�\EXCES���"R�QM�pb��� �R؋��"�QSCc �g��p�T_�p�X�`P9k�_�X/@K_��'R�v�HFB_8�FLI�C$Be�QUIRE�㱠�kO�k�zAuL< M^�� j �S��`_�u��2ef��MND�����P��������#sD����INAUT����֠I�=x N������	qQ�qPSTLb�� �4�LOCeRI�<�eEX�vANG�ڢQR�PODA�EŪ�P�*��MF Z�>��F�;"��E%����GFSUPN&� F�X�IGGW� � �s�;#��ܣ;# ��;$�R�X��h���w�X`L�SA�=QTII�� ��MFpn7B� t�pMDՁI�)�0 � A�qH�pX��DIA���ANSW������D�)taOR��2��P� `C�U �V,�O0�q�aOr��_2@��� �S0m�s4@��B����P��J�lЦ�P��KqE���!�-$B����}�ND2�2�1��2_TXD$XT�RA0�B��`L�OАP�
b1��r	L0��°f�Q�I��R�RR2�U� �0A���A�1 d�$CALI�P��G���2��@ ��!����<$R���SW0�4ݣCA;BC�xD_J��a\�p�_J3�
�G1SP�`\p�pP�B)�3(�k� �pX��JCh��2��O�I<¢qQCSKP�*��H���J�pRQ���ȵ��ȵ���p_AZ�2d���EL�c��1OCMP�sqQ0Q��cRThA%�C�1�e��1��1�G���U�Z�S�SMG��ƀDJ�Gb SCL�P�uS'PH__ pP�ų0z�p��RTERܠ�������_ q!`A�ЧpR��DI����23U��DF����LW��VE�L�!INP"��"�_BL0 �r*�â�1�x/�H�@�MECH��DTSA_ܡ�F�IN���A�P�f�H�Մ�q��� _wP ��մ����`��b%b�����.�DH�Pt���� $V��<s����$r��A�BV��$�1� RY���P�H �$B�EL��G��_ACCE0� \�Ak�OIRC_���c0�NT0Q�$PS�P�"L��p���# �Ё��q ���a���Dw���3��w��Q_�+����E[Pa�_M�G�CDD+��¡BFW� ǀg�G�w�b�<��DEe�PPABN6��RO��EE�# ��� ��#5A5`b�џ$USE_����P.G`CTR��Y��=�Z�1 ,�YN�PA��������M]Aq��B�%�O���"INC K��qd�K��RDá�QENC��L���r��Xb�T��IN�I�☋Ȁ��NT�A�N�T23_�¡B�L!OСB� �@I�`�t ��f�fPF�'e�GayC�РMOSI0��_b~���CpRPER�CH  g��A��  8�qC���D�� � ��������A��L��Zg���0��
���TRK��*!AYE��5a!��%#�p+�9aR1PMOM M��R5bf0k��tc�a"#���w�DU ��S_BCKLSH_C��%]@�@���PS�#k�*��CLALM�cAH �Ў�%CHK������GLRTY��������X1Ɓ_�_UMVCG6CVC9��_3�@7LMT%�_L)��x4��7E}=�0�;|0 ��5��:�\C��4|PCI|H3��`/��G5CMC!�9�=�C�N_��N �>Fp�S	FO�mV�򸁁��pA��EHCATN>SH���=�s81�!��B���B�H�,�PALN4B_PM51#_�����&,��#0T!5JaG�p`$S�OG1G>��TORQU��+� 
')s��b"��s�R_W`%$Q�,�T㨳U#�UI�[I�[I#�F�p�Qo�h~�5��VCa�0VaKe)b1�/n-�Co�5fJRK�/ltbgf_�DB��Mt��_�M:p_DL��GRV�T�d�d#�aH_H��c���j�COS�k-��hLN v`{2et�yr�y �QOz=|a�eZp"�aMYq�x�b�{��yTHET0�N�K23#��r�pC�B�vCB�C��AS����T����v�SB�.��uGTS����C,�
QK��C[�<d�Ls$DU0������1՘�@�Qx_��3�ANE����K .47������qA�u��p��e�h�aLPH�eׂ�ׂS2eJ�=uJ��Luׂ[vt�^�{v��V��V��3�VB�V�O�V]�Vk�Vy�V
��V��H�4�:�2���AQ�O�H]�Hk�H�y�H��H��O�OR�OƩ1�OB�OO�UO]�Ok�Oy�O��O{vFׂ�qY�=u^���SPBALANgCE_�q��LEE�H_�uSP��.v���=v��LvPFULC���ܲķܲLu��1��9�UTO_0!5Tg1T2�]�2N 1 h� =Ă�A!ް����X�\!T�O��j�P�INSEGh��R�EVb�� �DIF����1�����1���@OB���!�cn'2�P� 1�dLCHW3AR����AB Qp%�k�� �pm�b3X�!P�43������� 
4ҒQV�ROB,CR�v�(B���CT�_RT �� x $WEgIGH � $�d��3PI� IF��NE�LAG�2S܍�BIL��OD�J � ��STn���P���� ��:�@�џи£�
g T�Q  �2�	��DEBU���L�����MMY9���N�Cw�� g$D��S$a��.P�q ���DO_��A�ѹ �<��1�'�݁�B$���N���_�  ��O�  ��� %f0T� �e1Tx��Y��TICK����T1��%)� 2�!N,���,R� ���D���P���PRO�MPE� $IRuP'0����MAI�`L!��_�����! �R�`COD6�FU	 ��ID_K�������G_SUFF��P �����?�DOG���H���G�GR����$e�0�;��G�A$��@๺��H��_FI5��9�ORD� ��i�36�2���$ZDT����ྫ�4 *��L�_NA��2��D�DEF_I�j� P��C��C�<P�Jj�IS��v@��πC�D�P��Ag�4GA��2�D��"�6�D�rPO����LOCKE�AD�V�h��$ UM#�$<$ J$�0&#/0 Z0�&�;�Q ;�;<;�'�% ��P��s�Հ���W(5���TE|�!��( �џLOMB_2970���VIS�`ITY���A.QO�A_FcRI�a3��SI�c1��R/��7:��73O���Wf8Wr;�`h6rx`_�9EEAS�ӀE?Q`4�@���64�95�96��ORM_ULA_I�A�4wTHR�� �G�ѽ���p_�8o�COEFF_O�y��D$�M�G�A��S�Ј�#CAް���$ C����GR�� � �� $�P���X�TM�T��#, \��ER��T��n@�  �LLF:�S�_SV�rX�O@(5@༁paD@�{ �BSETUMEA�� !`���|��п � �@g� q�J@�Q܂�Q���V�2�����B�1Pcp��A��&k������REC��Q�S�K_���C� P~��1_USER9��)�xd���tx`9�VE�Lbx`���b�e��I�� ���MT��CF}Gna�  4�z��O"�NORE������b�OPWOR�ڀ �,��S�YSBU�aSOQPqd`bTzU{b��P��b9uPA{`��Q;s�aOP9 U���-q��3�p�mpI'MAG�PV�hp�3IMGp�uIN�0ar~�sRGOVRD��)s|`lqPnp�ss�πк ��u#�L�BT|΂�QPMC_E� qe�N�M�p�i�11n��qSLϰo`�� ���OVSL:b�S�"DEX�XP�����C_�ph�k  �ph�k r�����i⧃�Cd�� G������p_ZER�a/��Sna�� @ ҃=�O&��RI��M�
�� ����#2��E��o`�� H����ATsUS�P�C_T�qDXQ�B
P^�G��T�o�3�� o`� D ��jpS�Q���R���@Na�qXEX��U�������������W�U1Pd�yPX��~��g�g�3����P�G�e� p$SU�BF�=�g!F��JMPWAIT��w�^�WLOW"�F�M��#�RCVF��5�"Җa�RE��F���Cƹ�RL"�5�IG�NR_PL�DB�TB�P}#�BW����`U�थIG�Qqt�C�%�TNLNl�� �RT�sNO�0yNt�J�PEED��>Y�HADOW�!��`ERVEX�R�g��0�SPO� � L��:�r����CUN��!�~��RǐF��LY� _�P�,��PH_PKT�c���bRETRIEx��bnr  ɱv��FIҲ� ��мͰ�� 2��`D�BGLV��LOG�SIZ/�mRͰ~�U��7�D=��_TX�"�ME@CMa��EM�F�RW��"�CHEsCK�a�P�`�na� 0�鸌�A3LE	���PA���8bU��aPIP��na�� h $AR@*��� �W8�OH z�C@AT ��Wa*�`]���p�Ӥ�UX�`�͂ݑPL���d� �$�a�!SWITC�H"�WO����-�Y�LLB`���� $BAU`D�aBAM��0w�4�����J5n��a���6�ց�_KNO�W���ҿpUcADȢ��@}�D{`�PA�YLOA�Q� *�_P`�3�q3�Z0�Lg!yA�QHLCL_GP !�Pl��ѲaTy��r��F��CFPPg��Rj�u@Ig�RHP�g�!����B�0GP_�J����_Jq�aƐTAND��4b�hq��d��1PL��?AL_ �e�}��AbB�qF0CbD:/�Eb�J3$�8��� T��PDCK��p|aCO�P_AgLPHH��BE�P�H�Z���B��p� � �3�)�D�_10�2Z�D�PA�R������R�TIA46	56	6bMOM@BbOhb\�`Bu�ADBp�O�\PUBa�ARg�O���$0� 8���a��  E��M8�=��@T��kd�� e$PIF����a5�+��TO�+I7IEIS�������$�RO��,2��6�HIGt�6�v�o��o� v������#����<��v�SAMP�����:)�@#v���� o@n!GP��b}$�@�&o���) �bR� `;�%�1"�%IN�, �0##�(�+�$v��*8x�$;7;GAMM�%qSZ� �#�GET�CFI��Z���b
�A�IB�B�I����'$HI`�1A`��b�6E��8A�>�0�6LW�=�6�<�9F�6лB��:�CۥCH�K�p�`}�I_" бb�"��1�%��Gb�D��I8� ��$j� 1���@ItPRCH_D`�c"c���$`LE�a��a�X���@��M�SWFL���SCR	�100�r3�}$ �Q0�cU�'��B �)vY�o��UPI3AMETHO̓�Rۥ�R+AX)���X9��0N�ERI�T?$3k3IR���	���F�d$@!�# b�#b-iqL�@@!BeOOP�!p�QXa�!�QAPPQ"�F�p��\e}dhe�#RT�R7CO#�o�5E`�a��c�W�1�*a`����jS�bRA��kMG"���SVw�P0�CURHW�qGRO<� �S_�SA���t:u��NO��C�����:p�4�� ;�M�Y�z�{�,�xDOn�A�2i� ~%xZ�%������(�8�4��sp����X�M�
� � �CYQL)��'�QS��;>�Paa��C�����_�AC����M_Wip؂Hb�`փDfM��������7�AQT�PU�M+q�� ������YWJ�$�`L8� ]�J���H���H���H�\�ˠ�0N�Ќ3kӳSJ0X��O��1ZΕ���� ��bM�Cv|����@9 �aQ������_��� |{��:pb	�� O���:p;
����U
�zф5 h�w�r���^�x�P���P�MON_QUD  �� 8��QCO�U�A�QTHdpH�O��?�HYS�ES��?�UE*�0r��]O���  ڰP(���5[qRUN_TOⶃk��� P�&���CƁ��pIN�DE�TROGRA���OЗ�2H`NE_3NOӴ��IT�ְ�l�INFO��� �gѼ������E�O�I��� (�@SLEQ�'��'������OSZ@��� 4���ENABv���P�TION��ER�VE��ǚ�[�G�CFd�� @3�JX�1����0R����ϖǝ�_EDI�T��� �W�ݐK����1E�0NU���AUTVq�COPY��/ܚbp�M�1N9�=�RFPR�UT @�N��O;UC�$G���Ծ �RGADJ���[ h{�X_߀I�CP͐��ې��W��P�ؠP����Ч2N�_�CYCv�j�RG�NS`��x�BPLG�O_C�NYQ_FREQ�W"0�U�gSIZs�`@LA�S�L���]"0�CRE��0�S`@IFEǳNmAH!%��_G�SSTATU{��S~�MAILF"����P:�LAST���'��ELEMd�� �|apn�FEASIq� 8�s"lP_P��aCq>�b� �0IఔDL�0B��Ss�ABZ����Ḛ�V ��BA!S����2�U���Op$���RM� Rm�1 P��Ɠ��2��� F�)��惠	J� 2� �#���$0�� /��'�� ����[#TDOU���Dwb'��Pa �.�GRIyDڱZ�BARS�sTYrî�OTO������ y�_��!�����O̐a�� � ٰ�PORp����U�SRV���)DIXpT_��9K�U�U4�S5S6S7S8�7 �Fg2d��w�$VALU��-u0��o�i�F`��� !!m�c�ɱ���*x`AN,s���`Y�~.�TOTAL_��,q�;"PWB�I�P$REGENN*c"죁X����BE�&%�T1R����N!_S0p�'c  cV�����"��E��`D�-�%�#7V_H� DA%�� �0S_Y^qƒf�S�=�AR%�2� >��IG_SE;�� d��_���$C_��$CMr`k�|2DERmpD0�2IbAZ{3�U3v�ENHAN�C+�샠
m�8��i�1INT6����F���MASK�S��OVR�T�`pA�����OVC���
`��i¯O�|�+��PSLGM0>�� \ 6rg�_R)�8 ��Sł��1U^Q~��E�#�D�_U�DTE�� �O (�!�VJgF<Vrv�IL_Mu�&P1Vy�`�TQ%��S�߱��C����VS[CFa]P_%POpkSM�Y[V1�ZV1�[2�[U2�[3�[3�[4�[4�Zq\a�bpAcc�ǁ�IN,iVIB�5�[TH`�Od2Kh2�Wh3Kh3Wh4Kh4 Wh��jTw�fXplf`y'g$e8e$ePL��gTOR)�	�IN�ep	��@:r���d܀�MC_FH�]pB�Lqq�5. M�p1I�3;rw ��.���2܀KEEP_H/NADD4q!vt���yC���@�t�5r�@�sO�utC�3q+���s�7�sREM�r@�t����u�q�xU���e�tHPWD  ;vsSBM�1� ?COLLAB'��h�@,!���IT,�콐N�NO.�FCA9Lm�+#DON �A�r�� ,�FL|s���$SYN-p���M�Ch2�� U_P_DLY���w��DELAր����Y��AD%��� �Q�SKIPL�� Ą��O���B\R �P_�����������6� ��D���D�lC�yC� �C��C��C��C��9���RAa�� �XC0"�7MB�pN�FLIC����M�UxLz�GNO_H�x�rq��@SWIT��]Ր_PAͰGO� ��0�8U���W��V�F3�3NGRLTր���с �@�@8�3[���T_J��*��v�AP~0WEIG=H��J4CHq���cOR���BOO$ ��"]�~�J ���A0���5��OBY�Y��  �$�`AS=S�����A�F�MF� 6���S|��>�L�1b��$AAVM_W�RK 2 A���� 0  �#5H�������Ž ż	�ٽ���F�B���'��,� ؼK�W��]ϒϤϬ��p�BS���0 1�_�� < ������'�9�K�]� o߁ߓߥ߷������� ���#�5�G�Y�k�}� ������������� �1�C�U�g�y����� ����������	- ?Qcu����������C��A�XLMT\��n��  dIN#H5F@_ Fr�U�pC_O  �^�� ��
}I�D ?A�r ������(/ #/5/G/p/k/�M1�0����/zUPo@f��$  p�IOgCNVfBG �1P�&[�F�ǻ��� w 1}�P $m����]=a�Z?B�?� �&(}?�?�?�?�?�? �?�?OO1OCOUOgO yO�O�O�O�O�O�O�O 	__-_?_Q_c_u_�_ �_�_�_�_�_�_oo )o;oMo_oqo�o�o�o �o�o�o�o%7 I[m���� ����!�3�E�W� i�{�������ÏՏ� ����/�A�S�e�w� ��������џ���� �+�=�O�a�s����� ����ͯ߯���'� 9�K�]�o��������� ɿۿ����#�5�G� Y�k�}Ϗϡϳ����� ������1�C�U�g� yߋߝ߯��������߀	��-�?�Q�c�L�ARMRECOV� �,U64L�MDG �'�Q0�+��_IF F;6�/�"�4� F�T���w���������, 
�/��`�/ "4FT
$��x _�[�������'NGTOL  ��	 A  � >P{PPIN�FO �� ��������  ������/� 6/ /2/l/V/�/z/�/�/d����/?? (?:?L?^?p?�?�?�?��?�?PPLIC�ATION ?����� �HandlingTool E� 
V9.30�P/17_�7
�25793500�01,KV:CA-J1�09XAYN"O4B7�DF3(@�<CNo�ne�;FRA��? 1pM�6_�ACTIVEp� � �37  �CU_TOMODP���5�ECHGAPO�NL$_��;POUP�LED 1���� uPy_�_�_�KCUREQ 1	��W  T�Y�\�\	�_	e�0d���_�_ �_o"o4oFo�ojo����R��
E�dH�UxR�j?HTTHKY�o}o �o�o�o+=Oa s������� ��'�9�K�]�o��� ��폷�ɏۏ����� #�5�G�Y�k�}���� ��şן������1� C�U�g�y���寯��� ӯ���	��-�?�Q� c�u���Ύ���Ͽ� ���)�;�M�_�q� ���ϧϹ�������� �%�7�I�[�m���� �ߵ����������!� 3�E�W�i�{����� ����������/�A� S�e�w����������������UTO(_S�DO_CLEAN�E_�D|NM  - �_���� �^DSPDR3YR��EHI"P�@�~����� ��/ /2/D/V/�HMAX�0c��TW�t!XcsApRsA�BPLUGGcPdpSUWPRC5B� �m_/�"O�">P/SEGF<PK?,7 71��~?�?�?�?�?�/11LAP[n>�c O,O>OPObOtO�O�O��O�O�O�O�O7STO�TAL�&�)7SUSWENU[0h[ I�M_��PRGDIS�PMMC:0�!CLB1�!@@PhTOY�{&F5dS_STR�ING 1
4[
_�M-PS�J�
�Q_ITEM1�V  n�M�_o o%o7oIo[omoo�o �o�o�o�o�o�o!�3EI/O �SIGNAL�U�Tryout �Mode�UIn�p�pSimula�ted�QOut��|OVERR~X = 100�R�In cycl��u�QProg OAbor�s�Q�t�Status�S	�Heartbea�t�WMH Fa�ul��Aler (�XF�X�j�|�����p��ď֏� _ �[_�_�9�K�]�o� ��������ɟ۟��� �#�5�G�Y�k�}���WOR:0�[��)��� ݯ���%�7�I�[� m��������ǿٿ�p���!�3�PO�[ 	�Y�ͫB�|ώϠϲ� ����������0�B� T�f�xߊߜ߮�����T�DEV\���p��� $�6�H�Z�l�~��� ����������� �2��D�V�h�z�PALT���ͯ{������� ��#5GYk} ���������GRIy �[E�� m����� ��/!/3/E/W/i/@{/�/�/�/3+PR� �!]�/?#?5?G?Y? k?}?�?�?�?�?�?�?��?OO1OCOUO�/PREG���@?gO�O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_��_�_[}�$ARG�_��D ?	����<a�  	$[vW	[Ph]Pg�[w�qi/`SBN_CO�NFIGjp<k�q�r�a�aCII_SAVE  [t��a�c/`TCELL�SETUP �<j%  OME_�IO[}[|%MO�V_H�`	RE�P�,Z%jUTOB�ACK�a<i�b�FRA:\{Kc e{F�`'`�p9{G�x� �{�`� 21/�06/22 02�:23:42{F�rh{M�-�Z�Q��|��z�����ŏ׏���{F���)�;�M�_�q� �������˟ݟ�� ���7�I�[�m���� ���ǯٯ����!��� �  �q_}s_�\ATBCKCT�L.TMP DATE.D��h�z��������wsINI����u�fwsMESSAG�`ϱ�aD`�c�a�ODE_D�`�f�e��O���wsPA�USm� !�<k ,$	�r`x<eq��,		i� �ύ��ϱ�������!� �-�W�A�{�e߇߱��D�N�TSK  �Tͮ��zpUPDT��ͷd��XW?ZD_ENBʹ�j'�STA̵<a�.a�XIS�`UNT �2<e�a�`� �	 bf(� ��R��Lpv�+ ��jPg���	q  `	_�  �����p�����������5��� X�� 9�O >� i�� ?�k ���1���T���i�MET� 2���c� P��D{�%D���DJ��D���D���D?fa@����<䝲=T��<�z�=��=c�=u���6�.�p�SCRDCFG 1<e;�q ��e�bR�&8J\n� �{JZ���� %�I�{�{�@����<g�$}q�GRp��2�#C�N5A#p;k	}t&�_ED˰1��� 
 �%-I�EDT-�7z�/�/^� � u-}s|/{Jrbp�vu/^(?  ��52?�/k?�/O}��(G?�? �/?�?/?33�?6{ �?EO7��+O~O�?�?mO�?34�O&O_JO \N�OJ_�O�O9_�O35�_�O�__\N�_o ]_o_o�_36No�_ �o�_\Nwo�o)o;o�o_o37�og�o\N�C��o�+38�Z?3�~?��=�z� ��i��39��"���F���=ۏF�����5�Ï1CR?Uʟ ܟ�}���W�i������ X NO_DEL�/	"GE_UNU�SE/$IGAL�LOW 1;)�   (*S�YSTEM*A��	$SERV_G�RO"A�ʠN�REG�ӥ$��A�ʠNU�M����PMU|v�A�LAY���A�PMPA�L�Q�CYC10�W�j�T�X���UL�SUJ��l�N�գ�L��ߴBOXOR=I��CUR_̰��PMCNVF��̰10��2�T4�DLI2�ſ�	*�PROGRAҤ?PG_MIX���F��ALbšϋ����B��ʮ$FLU?I_RESUp�����.�MR��(�(�9�r߄ߖߨߺ� ��������&�8�J� \�n��������� �����"�4�F�X�j��|���i�LAL_OUT ���#*!WD_ABOR� �����ITR_RT/N  �$�")��?NONSTOO � ��CE_RIgA_I��c �&!M FCFG �;*cZl_�PA��GP 1.v����x��CH  #Up%�%�%�%��%�%�  DV��DQQ QӠD4Q>Q$��%x�E�%�VQ	�Z"�/QY;�$DT�aQ�m�zQ�@ Dˉ��&?�M HEE�ONFI:�����G_P�1v b�;%///A/S/�e/w/�/�/�KPA�US�1 %c� ��$�	��=���n>������	�,�$?��z�?ј���N��??�u? C?)?g?y?_?�?�?�?��?�?�?	O�?-O�.M~ NFO 1 %��  � �	��O �p@� 9�W�n`�����B�[MBXz�^��VxĴ��&� D�L��Ī-�C~���@�Q�A�߶B:�J�A�������/D`���A<sA�*I�9�M O�pv��ALL�ECT_p^F��WENb���:R�ANDE&S�.W��#�1234567890�W��䡆�_�V�
 p�� �)�_�_��_ �_Co�/ o2o�oVoho zo�o�o�o�o�o�o 
c.@R�v� �����;���`*�����jT�2.[� X=[lRIO # wY:Q����%�7�χTR� 2%!��(� �
`�E���"ލo��BV_WMOR��#� < .���oA������4�"�X�F�ђ���$
ߝ,�?��@��R� K��^�P�B	&._����%��Y�
�W�W��}��@���Ea���� �sj�AVP�DBϠ(��n�c?pmidbg����L �:�d��p�|B��  �d�翆�Q�Le�0�l��R����mg�����e�f�`�!Me�>r�ud1:�߮����ǱDEF '�H�)��c��b?uf.txt���\��Ű_MCؓ)�����dL�-�ה*;�x�z�]=4�#�Bpp@B�B<B��g+B���B���B��PB��IC�ۿ�I�CZ��C����C���C�'��C�X�C���E�k�IE�>�\E��KE��FE�k#E����E�o�F�١\�l�-⁧,���W �
H��P��Z��l����x����%hCdO7������.f�[rٚExD��l�E�G([����*f�E-x� F��t�fEпU�H�i���  >�33%�>���?����n����5ِ���H���A����L_��<#���������C"H%�RSMOFST %�ڼ=OKFP_T1��-Ƴ�A`ť�MO�DE .ӯ���x� �A;�6�XR?��<�M�>���%�TES�T��+���R(R/�_�~�x�A����T�@k�$C��B�������C��@����@:d��� 4�oA�
/�*gIpS0q?&#���1ߝ�TW�RT_~��PROG ��y%�/d׀NU?SER  WU�!��Rh#KEY_TBOL  ߕ�!iB��	
�� �!"#$%&'()*+,-./�W�:;<=>?@A�BC��GHIJK�LMNOPQRS�TUVWXYZ[�\]^_`abc�defghijk�lmnopqrs�tuvwxyz{�|}~��������������������������������������������������������������������������q1���͓���������������������������������耇�����������������������k LCK�,y�$�� STAT�?e_AUTO_DOTV9x/CINDOTNbQR�:O,FT2xO��%STO�P_O�@T{RLm LETETW��J_SCREE�N ߚk�cscERU�@MM�ENU 12λ <�,�/M_�%,_ V_�_u�h_�_�_�_�_ �_�_�_3o
ooBo{o Rodo�o�o�o�o�o�o �o/e<N� r������� �O�&�8�^���n��� ͏�����ڏ��K� "�4���X�j������� Ɵ��֟�5���k� B�T�z���������� ү����.�g�>�P� ��t���ӿ���������Q�o�S_MA�NUAL�O�BZC�D,"3�	�"�"��L��?|(��L��5�4�Bȁ��#��DB;COV@RIG�GI���_ERRLs 	5;�(�ςߔߦ�� /�NUMLI�M�CT�y% DB�PXWORK 16;�q���*�<�|N�-DBTB_�AG 7^ݕ����DB_AWA�Y7�(GCP ry=��_AL��O��3�Y�@�EyjFܤ�Q� 18� , 
��_!^���^�X!�^�h�_MU@I� ��@% x�ONTImM�G�y������
�%�MOTN�END�/�REC�ORD 2>^�� �f�g�G�O� .g���Zl~� '��.�R +��a���� ���z/r'/� K/]/o/�/��//�/ 8/�/�/?#?�/G?�/ k?�/�?�?�?�?4?�? X?�?|?1OCOUOgO�? �O�?�OO�O�O�O	_ xO-__&_c_�O�_�_ �__�_�_P_ot_)o ;oMo�_\o�o�_�oo �o�o�o�o�o%�oI �om��>�6 �Z���,�>��q��TOLERENC��B����L���/�CSS_CNS�TCY 2?�����H���谏��Џ �����*�@�N�`� r���������Пޟ�����DEVICEw 2@�� �� R�g�y���������ӯ����	�g���HND�GD A����C�z���LS 2B<����������ӿ�������PARAM C��d�d�y�~\�RBT 2E�ۗ8L�<Y��� C������  É��������Ɗ��ǂ��Hl����\���@�����C�˭Ó��� B7�  ��<�O��%ӓ�&�C�]�D#� ����4B۠�Y�^Ԡ���	�c6� ��	�I��ߞ߰����� ����E��.�{�R�d�|v�	�C�$�DN��D���� 	 �B!ffA����A_33A1�w�AU�����	�����B�|�����C����^��B+B.2�q33�Br2������P�b�.��33 �X� `� ����g��	�qÓ�� �����������P '9�]o��� ���:#5 GYk���� / {�/*//N/9/r/]/ �/�/�/�/����? �/�/J?!?3?�?W?i? {?�?�?�?�?�?�?4O OO/O|OSOeO�O�O �O�O�O�O�O0_�/T_ ?_x_�_u_�_�_�_�_ �_�/�/_�_�O'o9o �o]ooo�o�o�o�o�o �o�o:#pGY k}�����$� ���l��_��{��� ��؏�Տ���2�o ;�M�z�5�c�u����� ����ϟ�.���)� ;�M�_�������⯹� ˯ݯ���`�7�I� ����#�̿���ۿ� ��8�J�5�n�I�w��� �ύϟ���������4� ��j�A�Sߠ�w߉� ���߿�������T� +�=�O��s����M� �����,��P�;�t� _������ϳ������� ��(��#5GY �}������ �Z1C�gy ����/��2// //h/S/�/w/�/�/�/ �/���/�??d? ;?M?�?q?�?�?�?�? �?O�?ONO%O7OIO [OmOO�O�O�O_�O �O�OJ_�/n_Y_�_}_��_�_�_�_�_oZ��$DCSS_SL�AVE F����?a�~(j_4D  ?n�TcAR_MENU G?k o�o�o �o�o�o�o&R�o$�6$nuaSHOW �2H?k �  .R#Q}�u�o�������*�<�N�  vp��������͏ߏ ���'�9�`�Z��� ��������ɟ۟��� �#�J�D�n�k�}��� ����ů�����4� .�X�U�g�y������� ֯ӿ�����B�?� Q�c�uχϙ������� ����,�)�;�M�_� q߃ߪ�$߹������ ��%�7�I�[�m�� �ߣ������ ���� !�3�E�W�i������ ���������/ ASz�w����� ����+=d as������ �//'/NK/]/o/ ��/��/�/�/�/�/ ?8/5?G?Y?�/z?�/ �?�?�?�?�?�?"?O 1OCOj?dO�?�O�O�O �O�O�OO�O_-_TO N_xOu_�_�_�_�_�_��Op_ooICFG7 I_eiciQ�PqdMC:\�WpL%04d.C�SV$ofPcpoPr��PqA �cCH�`z@HV�o?_�o�oiQ��V��bq y�ajpGJP�2s�n�afP�G}6dRC_OUoT JBeLa�Yr)o_C_FS�I ?y D{�V��� ���+�T�O�a�s� ���������ߏ�� ,�'�9�K�t�o����� ����ɟ۟����#� L�G�Y�k��������� ܯׯ���$��1�C� l�g�y���������ӿ ����	��D�?�Q�c� �χϙϫ��������� ��)�;�d�_�q߃� �ߧ߹��������� <�7�I�[����� ����������!�3� \�W�i�{��������� ������4/AS |w������ +TOas �������/ ,/'/9/K/t/o/�/�/ �/�/�/�/?�/?#? L?G?Y?k?�?�?�?�? �?�?�?�?$OO1OCO lOgOyO�O�O�O�O�O �O�O	__D_?_Q_c_ �_�_�_�_�_�_�_�_ oo)o;odo_oqo�o �o�o�o�o�o�o <7I[��� ������!�3� \�W�i�{�������Ï �����4�/�A�S� |�w�����ğ��џ� ���+�T�O�a�s� ���������߯�� ,�'�9�K�t�o����� ����ɿۿ����#� L�G�Y�kϔϏϡϳ� ��������$��1�C� l�g�yߋߴ߯����� ����	��D�?�Q�c� ������������� ��)�;�d�_�q��� ������������ <7I[��������!��$DCS_C_F�SO ?����M P '!j�� ������#// 0/B/k/f/x/�/�/�/ �/�/�/�/??C?>? P?b?�?�?�?�?�?�? �?�?OO(O:OcO^O pO�O�O�O�O�O�O�O  __;_6_H_Z_�_~_ �_�_�_�_�_�_oo  o2o[oVohozo�o�o �o�o�o�o�o
3. @R{v���� �����*�S�N��`�r�������3C_RPIJ\��� 0�+�֏I��<�����,��6SL�@z��� �.�)�;�M�v�q��� ������˯ݯ��� %�N�I�[�m������� ��޿ٿ���&�!�3� E�n�i�{ύ϶ϱ��� ��������F�A�S� eߎ߉ߛ߭������� ����+�=�f�a�s� ������������ �>�9�K�]������� ������ԟg�����# LGYk���� ����$1C lgy����� ��	//D/?/Q/c/ �/�/�/�/�/�/�/�/ ??)?;?d?_?q?�? �?�?�?�?�?�?OO <O7OIO[O�OO�O�O �O�O�O�O__!_3_ \_W_i_{_�_�_�_�_��_�_T�NOCOD�E Kk���U�PRE_C�HK Mk��PA� �P�<� �`k�so�ok� 	 <go�o�o�o �o�o'9%o �[������ �#�5��Y�k�E��� ���o��׏鏃��� ��+�U�/�A�����w� ��ӟ��ߟ	����?� Q�+�u���a������� ŏ�����;��'� q���]�������ſ� ɿۿ%�7��[�m�G� yϣ�}Ϗ�������� !�ۯ	�W�i�Cߍߟ� y����߯������� A�S�-�w��c�u�� ��������+�=�3� %�s������������ ������'9]o I{����� #�/YO�a�� �;����// �C/U///a/�/e/w/ �/�/�/�/	?�/??? ?+?u?�?a?�?�?w �?�?O�?)O;OO_O qOKO]O�O�O�O�O�O �O_%_�O_[_m_G_ �_�_}_�_�_�?�_o !o�_EoWo1oco�ogo yo�o�o�o�o�o A-w�c�� ����_�_+�=�� I�s�M�_�������ߏ �ˏ��'���]�o� I��������۟��ǟ �#���G�Y��A��� ��{�ůׯ������ ��C�U�/�y���e��� ��������	��-�?� �c�u�k�]ϫϽ�W� ��������)���_� q�Kߕߧ߁߳��߷� ���%���I�[�5�g� ��ϙ�����s���� ����E�W�1�{���g� ������������/ AMwQc�� ������+= asM����� ��/'//K/]/7/ I/�/�//�/�/�/�/ ?�/G?Y?�/}?�? i?�?�?�?�?�?O�? 1OCOOOOyOSOeO�O �O�O�O�O�O_-_#? 5?c_u__�_�_�_�_ �_�_�_o)oo5o_o 9oKo�o�o�o�o�o�o �o�o�oI[5 �K_y����� �3�E��1�{���g� ��Ï�����ӏ�/� A��e�w�Q������ ��������+��7� a�;�M�������ͯ߯ ������K�]�7� ����m���ɿ��џ�� ϫ��G�!�3�}Ϗ� iϳ��ϟ��������� 1�C��g�y�S߅߯� �ߛ��������-�� �c�u�O������ ������)��M�_� 9�����o��������� ��7I?�1 �+������ �3Ei{U� ������/// 	/;/e/[m�/�/G/ �/�/�/�/?+??O? a?;?m?�?q?�?�?�? �?OO�?!OKO%O7O �O�OmO�O�O�/�O�O _�O5_G_!_k_}_W_ i_�_�_�_�_�_�_o 1ooogoyoSo�o�o �o�o�o�O�o-�o Qc=o�s�� �����#�M�'� 9�����o���ˏ��׏ ��o	7�I��U�� Y�k���ǟ�����ן 	�3���i�{�U��� ���������ӯ�/�����$DCS_�SGN N��[����t��22-DEC-2�2 00:17 ��d�JUN-21? 02:29u������ T�@�R��R�S��������`�4�����Þ諷�ì�  G�V�ERSION �S�V4.2�.14ݻEFLO�GIC 1O���  	���$�7�$�F���PROG_ENB  ��.Ñ�g�ULSE  L����_ACCL{IM���������WRSTJN�T��[��C�EM�Op̐������IN�IT P&�����OPT_SL �?	���
 	�R575��Q�7�4V�6W�7W�50
{�1{�2W�8ȥ��>4�TO  @ݯ�t���V�DEX���d[����PAT�H AS�A\TINKER\ ��f�x��HCP_CLNTID ?��.� 8Ȱ�����IAG_GRP� 2U�_ ���"'��FCP FV�� ��Ez 	�@<����B�  &����#�,�O�=�Cp � C��C��� Ck�Cn.ߘCb���mp5m8 78�90123456�����'��  �A�(�A�����  AͮA���A�ffA��\)A���\�A��װ�����@)���u�Aw�A��+�SA�,���Bu�BɎ�� ��@؎�
���B5=qB0f�fB+p�B&Q��B!
=B��B�B` 	h z����	��/ �C	&z��B"` � ���Bh h 	�R�BQ�A������v����D�AH��AC��=�A8��2=q�A,��%�A/�Ah �$6HZX��A_S
=AM��G�}@h:{A3���,� $��AG�������\Z���Tz�AN��H�� B ;��4h-A& ff /,/>/P/b/D3�? �?M?_?�/3?}?�? �?�?�?g?y?�?%O7O@O[OmO�?yO$����^� v!� �=�G�=u�A>�Ĝ�E�7'���7� P{��6�7�
U�@ʏ�\&V�p�2U��@f Ah��=PA� ��<N�W;�
��<�%�=�U*�=��k=�@�^�;'�U<�X�����>��C�  <(�U.�� 4"R�� �U�����U��A�? ��Oo�MoDoVo� �Tbo�o&o�o�o�o�o��o�I?S��?H��9?,I�?&��y&u���@BG	���� S��"wt
�x,�,�!�p�r�33f�x��������|�p���"3���~E�@ E�� Z�D+�f����� ���P���ÏՏ��� �{�$��{B�H����D�L�Ī.�C~�H@�V�A�:B:� T������������˟���=�����=R
�=��^��M����d6
_Q�P�B8?Q�;ě�^����CT_CONFI/G V���Ò��egM���STBF_TTS�ǁ
ɮ�Ó����G�MAU��t��M_SW_CF��W���  ��G�OCVI�EWՠX�!����g�y��������� ��U����� �2�D� ӿh�zόϞϰ���Q� ����
��.�@�R��� v߈ߚ߬߾���_��� ��*�<�N���r�� ��������m��� &�8�J�\���������������j�RC�Y�e�!v�܎G6�kZ�~�ǤSB�L_FAULT �Z
*��GPM�SK���2�TBRF�[�L��� ��(Tf��TDIAR\��!���[Q�UD1: �67890123�45���[Q���P 6�//)/;/M/_/ q/�/�/�/�/�/�/�/@??�v�9�R
�<[?�RECP��
��?��;��?�? OO&O8OJO\OnO�O �O�O�O�O�O�O�O%?�7?I?F_+�UMP_?OPTION����`QT���	�UP�ME��t_Y_TE�MP  È�k3Bg��P�Ag��TUNI󠹥�Q��YN_BRK �]@�+�EDITO�RfQlQ�_#b_x0E_NT 1^	4�,&
ROS_W�ILD;�LL A�VE H w`AM�|aZ&AVIZ�MOu`oo�k&�NORM_TO_�DRI�o�kTO�OL_1_PICOK_LE�o�h�i?APROAC�o�d��b2�`OPOF�F�f-&PL�CHANDSHA�KE OW&B|"u��e2�o�t��t"�jSCI_�TAIL_SWI�T� ��dPF�c�PCLA�Q0��d�J�U�Z�T&�AU�`CALIB8�d��S4&fa�a�SMie����&
>M�20_3 ��ޏ>l�WRITEnp���
��fTRANS�PORT_POSy �F�SAFE[��IiR`��h�a��Z�E���`���"`MGDI_STA�U�J��Q�� "`NC_INFO 1_�5R���L�����(���ܒ1`� ��_i�\�v�
v�d 6_ïկ�����/� A�S�e�w��������� ѿ�����+�=ώU T�f�xϊϘɰ��Ͼ� ��������*�<�N� `�r߄ߖߨߺ����� ����&��M�W�i� {��ϱ��������� ��/�A�S�e�w��� ������������ +E�Oas��� ����'9 K]o����� ���/#/=+/Y/ k/}/��/�/�/�/�/ �/??1?C?U?g?y? �?�?�?�?�?�?�?	O O5/G/QOcOuO+O�/ �O�O�O�O�O__)_ ;_M___q_�_�_�_�_ �_�_�_oo-O?OIo [omoo�O�o�o�o�o �o�o!3EWi {������� ��7oA�S�e�w��o ������я����� +�=�O�a�s������� ��͟ߟ���/�9� K�]�o���{�����ɯ ۯ����#�5�G�Y� k�}�������ſ׿� ���'��C�U�gρ� ���ϯ���������	� �-�?�Q�c�u߇ߙ� �߽���������1� ;�M�_�q�ϕ��� ��������%�7�I� [�m������������ ����w�)�3EWi �������� /ASew� ������/! +/=/O/a/{�/�/�/ �/�/�/�/??'?9? K?]?o?�?�?�?�?�? �?�?�?/O5OGOYO s/iO�O�O�O�O�O�O �O__1_C_U_g_y_ �_�_�_�_�_�_�_O #O-o?oQoo}O�o�o �o�o�o�o�o) ;M_q���� ���	oo%�7�I� [�uo�������Ǐُ ����!�3�E�W�i� {�������ß՟��� ��/�A�S�m�w��� ������ѯ����� +�=�O�a�s������� ��Ϳ߿���'�9� K�e�WρϓϥϷ��� �������#�5�G�Y� k�}ߏߡ߳������� ����1�C�]�o�y� ������������	� �-�?�Q�c�u����� �����������) ;Mg�q���� ���%7I [m����� S/!/3/E/_i/ {/�/�/�/�/�/�/�/ ??/?A?S?e?w?�? �?�?�?�?�?�OO +O=OW/aOsO�O�O�O �O�O�O�O__'_9_ K_]_o_�_�_�_�_�_ �_�?�_o#o5oOOEo ko}o�o�o�o�o�o�o �o1CUgy ������_�_	� �-��Yoc�u����� ����Ϗ����)� ;�M�_�q��������� ˟����%�7�Q� [�m��������ǯٯ ����!�3�E�W�i� {�������ÿտ��� ��/�I�S�e�wω� �ϭϿ��������� +�=�O�a�s߅ߗߩ� ���������'�A� 3�]�o������� �������#�5�G�Y� k�}������������� ��9�K�Ugy �������	 -?Qcu�� �������//)/ CM/_/q/�/�/�/�/ �/�/�/??%?7?I? [?m??�?�?�?//� �?�?O!O;/EOWOiO {O�O�O�O�O�O�O�O __/_A_S_e_w_�_ �_�_�_�?�_�_oo 3O=oOoaoso�o�o�o �o�o�o�o'9 K]o�����_ ����+o!�G�Y� k�}�������ŏ׏� ����1�C�U�g�y��������� �$E�NETMODE �1a,���  �p�p��u���ؐOATC�FG b,���?��C��$�DATA 1c��A���*w�*�������˯ګdگ��0��v��)� ;�M�_�q������!� ˿ݿ���%ϟ�L� ÿm�ϑϣϵ���A� S����!�3�E�W�i� ���ϟ߱��������� s� ��A�S�e�w�� ���'����������+�=�ؐRPOST�_LO.�e`���
�E��������בRR�OR_PR[�%��%������TAB_LE  �6��:L^G�RSEV�_NUM ��  � Q��_AUTO_EN�B  ����_;NO� f��}�  *�� ��� �� �� � +�� �#�FLT9R��HIS����퐸_ALM 1]g� �����p+$�����//(_��   ����^*ؐT�CP_VER �!�!��)/$EX�TZ�_REQ_9�	�#SIZ�/�$�STK�)��~�"TOL  ��{Dzg�A �$_BWD> 0C?1��(3DI-1 h�2�j�	���D;STE�PU?g?ؐ�0OP_�DO�/֑FACTORY_TUN_�d�9DR_GRP� 1i�Id 	�Y/O�@��������6��Mj�����~ ��� ���OBC]OnM XO�O|O�O�O�O�O�O �O�O3__W_B_{_�
 K1���_�_W$__q_�_�_o��WC��NC� � C�  B��yh;e�]@UUUWo�UU�_�oo E׻� �o��^P]���P�W�Pm�4�M�D�aL��om?�`�o�o�:N�:�o�:I��9-��+uon$��������1�T��KG�F���ЗFE�ATURE j�,�?0�H�andlingT�ool �u���English �Dictiona�ry�w4D St΋pard�v�uAn�alog I/O��w�wgle Sh�ift�uto �Software Update��matic Ba�ckup�y<�gr�ound Edi�t�p�wCamer�a�pF�CnrR�ndImA�x�om�mon caliOb UIs���nZ����Monitor���tr�pReli�ab�p�xDHCP����ata Ac�quis�ia�gnos8��q�i�splay]�Li�cens��oc�ument Vi�ewe΂�ual� Check S�afety���vhanced���z���ss�Frk��wxt�. DIO ��f�i;�ϗend��E�rr̀L:��×s��r�pڐ .0�zF�CTN Menu�v�=�TP I�n,�facS��uG�igEe�w�S�p �Mask Excڠ�g̗HTc�Pr?oxy Svt���igh-Spe���Ski��˥3�ސm�munic7�ons�urJ�,� ��q�f�connect� 2�ncre�sGtru�r�C�ej��J:�ˤKARE�L Cmd. L橠ua��z�Runw-TiːEnvp�^-�el +;�s9�S/W�wU���s���Book(Sys�tem)�zMAC�ROs,ܢ/Of'fse���Hސ!�����MRǀÂ9�MechStop��t3����i�� �o�ax���p9�.�od�pwitch��C�.�y.$���Optm�ϜCû�fils�B�g����ulti-T���]��yPCM funM�K�o���D�^k�Regi��r �N�ril�F[ۣ��pNum Selg�|��ɐ Adju����� ���tatu���n��uRDM �Robot�pscgove�qK�ea<��ːFreq An;ly �Reme�ޑ�n�wK�W�Serv�oސ���xSNPX� b���SNc�C�lik����Libr�s��p v� ���oٰtJ�ssagD�ˤr  ���{r �/Id�G�MILI�Bp�J�P Fir�m�Z�PJ�Acc<T�\�TPTX��H�eln���K�q��[�orqu�pimGuláq�u���Pa��Z�S����&κ�ev.G��ri�����USB poort ��iP���al��R EVN�T�� nexcept����yԗĘ���VC��r���k�V@���) �#S��sSC��[SGEp�fUI�{Web Pl&����� ���j�!�ZDT A�ppl���z
!EOATV�@��v��A'Grid[�M�;-//iR.�z�&.��0N�-2000i�C/210L�|2D Gui� m����wGraphicܽ�uDV-��Pa?th Ctr�s;�ף.5�udv��DC�SO ck���ula�rm CauseM/��ed�x�S�p�8 rityAvo�idM��l�pāGAu�v�?�2g1��s�pt(3x�yc�p������ ���d1os./ףc��H���r/���trans.be�tw.V�_�mai�n Nʑ��.w�a�n.����Axi1sޑ݁?�RAO ɐ`�;�,����/C��oq����*1������8��h4�zNRT^�%�On�pe Hel���O�ROFINE�T CP16XX FW�@O՝Кр!�tr�ROS Eth�Cg1e '�������7 �2���	2��s�*sup�t̓p!�iR*� Pk�jfGiG԰k�cm�Im��F�k�nn�sp3�va�$64M?B DRAMw_�c�FRO�o��<�x���a�ell�|��shKqWiwc��fu�YpQ{|ty�ps������r��%^Cr��� �BO�`*A��{���E��MAIL���t@@���뗝V���q���T1ǀ��KףƷn�ear[� m���R��*\0pŃ��o�Qb�o�1dri��UP#T c��O��c:���g�4pk Syn.�(RSS)g�quir �O�.W� ��$8��ϰ��uesjE�UCma׺��`����S-@duk ��p��smi�)3DL&�M��a���d"K��l� Bui<�n�A'PLCh���VQu�sCG��߯CRG��b�DW��#�LS,�&�BUH��Kñg�&iTA����B���qU��TCBԿ涛�巋�F(��ׯ�pG�����TEH������V�Ϫ�o�!F���ӿ�G�Qא?�Q�{��H���IaA���֯��LN����Mw��_����	N���P�߅�[��	R#��S��������W���s��VGF7�I�P2+�e��e�$S�e�D��e�FC�e����,TUT��01���2TBG�G��;ru@�0 U9I��%HMIm�ponT��'HDfor �b���f�C�f�BI/��mTPG����F SWIME�ST�V257935�$��"&/ \Se����� ���"//+/X/O/ a/�/�/�/�/�/�/�/ �/??'?T?K?]?�? �?�?�?�?�?�?�?O O#OPOGOYO�O}O�O �O�O�O�O�O___ L_C_U_�_y_�_�_�_ �_�_�_o	ooHo?o Qo~ouo�o�o�o�o�o �oD;Mz q������
� ��@�7�I�v�m�� ����ЏǏُ���� <�3�E�r�i�{����� ̟ß՟����8�/� A�n�e�w�����ȯ�� ѯ�����4�+�=�j� a�s�����Ŀ��Ϳ�� ��0�'�9�f�]�o� �ϓ��Ϸ��������� ,�#�5�b�Y�k�}ߏ� �߳���������(�� 1�^�U�g�y���� ��������$��-�Z� Q�c�u����������� ���� )VM_ q������� %RI[m ������// !/N/E/W/i/{/�/�/ �/�/�/�/???J? A?S?e?w?�?�?�?�? �?�?OOOFO=OOO aOsO�O�O�O�O�O�O ___B_9_K_]_o_ �_�_�_�_�_�_o�_ o>o5oGoYoko�o�o �o�o�o�o�o: 1CUg���� �� ��	�6�-�?� Q�c�������Ə��Ϗ ����2�)�;�M�_� ��������˟��� �.�%�7�I�[���� ������ǯ�����*� !�3�E�W���{����� ��ÿ����&��/� A�Sπ�wω϶ϭϿ� ������"��+�=�O� |�s߅߲ߩ߻����� ����'�9�K�x�o� ��������������#�5�G�t�  � H552�f��21��R78���50��J614ޒ�ATUP��54�5��6��VCAM��CRI��UIFv��28��NRE���52��R63��S�CH��LIC!DwOCVRCSU���869��0��EI�OC"4��R69���ESET����J�7��R68��MA{SK��PRXY
]7��OCO�3��h��� ��3�J6���53uH'LCH^�OPLG��0�MHCR�SpMkCS��0�55���MDSW�OP�MPR6 50n��PCM	R0 '�� ��z551��5u11(0��PRS��69�FRD��FwREQ��MCN��{93��SNBA.^(SHLB�&M�'t6 �2��HTC���TMIL��uTP�A�TPTX�&EL�&zu8�����wJ95TUT�95�UEV�U�EC�UFR��V�CC�8O�VIP��&CSC!6CSGt!g I��WEB��7HTT��R6,C8l���6CG�7IG�7oIPGS*FRC�&�DGH7�R9nT'R76��R8��@qG85uR66�qG51�53%'6�8}G6626�1(6J74��7Y5�H�H51R?�R5\76 9Rk58aW88854eGq6|G
P��NVD��R6|R77}G7�9�4W87aW68qGk(R7� �D0|GFhRTS�&SVMCLI���CMS�f`���STY�'6�CT�O��f �7tNNvWNN�ORS�� ��EXTAF6 }X_(6 �OB�I�h�WR67uCPR��'L�7S�j1��6�7�SVSESL�M�V3D�8P�BV!6APL�A�PVEgCG��CC�RqCD�7CDL�AFCSBiCSKv�CT7CTBGTB�7TC�&F�%�`PF�	F�EgTC�;TC�CTEE����wTE]���7TF*1�F=�G%�Gى���H��I�&���,7C�TM=�DhTM�N*��P�P%�R1�hh�TS1�W��AFVGmF��P2�7P2�&TƐ��D��F	V'x�VT�����VTBZ�wVhIH�'VJ@n��KLVigVK�7=V�7Gene��m� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t����������� ��(�:�L�^�p��� ������������  $6HZl~�� ����� 2 DVhz���� ���
//./@/R/ d/v/�/�/�/�/�/�/ �/??*?<?N?`?r? �?�?�?�?�?�?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb�ty  H�55�pq�q��sR�78�|50�yJ6;14�yATUq��t�545�|6�yVC�Aɔ�sCRI�U�Im��u28�NR�E�z52�R63�{SC���sLIC^U�DOCV��C4���t869�{0�zE�IOM�\�4�zR6=9�ESET�{��J7�R68�zM�ASK�yPRXY�6�7�zOCO�3��|�z"��|3u�J6��|53ŊH��LC�HU�OPL)��u0^��MHCRV�S��MCS�|0%�55��zMDSWv���OP��MPR��r�Ŝ�0�zPCM5�R0`ԫ"��z"�ś51�{�51�0�zPRSv�69u�FRD%��FREQ�zMCN��z93�zSNBA�f���SHLB��M�Իr�e�2�zHTC��zTMIL�|ŊT{PA�TPTX�#EL��"�ŋ8�{�p�u�J95E�TUTv��95u�UEV�wUECU�UFR%��VCC��O5�VI�P%�CSCU�CS�GU���I�yWEBn�zHTT�zR6d�؃��pU�CGt�IG�T�IPGS��RC�%�DG��H7t�R�9D�R76�zR8�d�2��85ŊR6m6�51��53�[68%�66��2��u6�6E�J74�{�75E��51E�RFӜR5��r���9���R58U�8t�54��6$����zNVDv�R6$�R77%�k79��4��87U�368�c�R7D�B��E�D0$�FSRT�S��SVM��CL9I���{CMS劲 ��zSTY%�6t�C�TO�z���7ČN�N��NNu�ORS85�B��zEXT��r��%�S�r�u�OB��I�e��R67ŊCPUR��L�SC1u��67u�SVS��S;LM�V3D%�4�wPBVU�APL劷APV�CG�zC�CR�CD�CD�L��CSB��CS�K��CTD�CTB6��TB%�TCպ20�<��205�20�TCv�+TC�CTE����0�+TE���05�TUF<F%<G<G�=
�<H�<I��B@�<d�gCTM%<�TM�,UN�<PELP<R<��TS<W�M��V�GF[P2��P2���2P%\D%\F5�VƳVT�{�P��VT�B�+V��IH�V��ЖyKLV�VKz%�Vt�Gene�x ux,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� �,�>�P�b�t����� ����������( :L^p���� ��� $6H Zl~����� ��/ /2/D/V/h/ z/�/�/�/�/�/�/�/ 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4oFoXo jo|o�o�o�o�o�o�o �o0BTfuu}~pSTDyt?LANG�t�y �������+� =�O�a�s��������� ͏ߏ���'�9�K� ]�o���������ɟ۟ ����#�5�G�Y�k� }�������ůׯ��� ��1�C�U�g�y��� ������ӿ���	�ϸ-�?�Q�RBT�vOPTNnπϒϤ϶� ���������"�4�F� X�j�|ߎߠ߲�����8�����DPN�t$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������//�&/8/J/\/�uted �tqx�/�/�/�/�/ �/�/
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__ &_8_J_\_n_�_�_�_ �_�_�_�_�_o"o4o FoXojo|o�o�o�o�o �o�o�o0BT fx������ ���,�>�P�b�t� ��������Ώ���� �(�:�L�^�p����� ����ʟܟ� ��$� 6�H�Z�l�~������� Ưد���� �2�D� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬϾ������� ��*�<�N�`�r߄� �ߨߺ��������� &�8�J�\�n���� ���������������(�:�L�^�p�99�r��$FEAT_�ADD ?	��������  	q��������� ��0BTfx ������� ,>Pbt�� �����//(/ :/L/^/p/�/�/�/�/ �/�/�/ ??$?6?H? Z?l?~?�?�?�?�?�? �?�?O O2ODOVOhO zO�O�O�O�O�O�O�O 
__._@_R_d_v_�_ �_�_�_�_�_�_oo *o<oNo`oro�o�o�o �o�o�o�o&8 J\n����� ����"�4�F�X� j�|�������ď֏� ����0�B�T�f�x� ��������ҟ���� �,�>�P�b�t����� ����ί����(��:�L�^�p�������D�EMO j��   q�۽ѿ ����F�=�O�|� sυϟϩ�������� ��B�9�K�x�o߁� �ߥ����������� >�5�G�t�k�}��� ����������:�1� C�p�g�y��������� �� ��	6-?l cu������ �2);h_q �������/ ./%/7/d/[/m/�/�/ �/�/�/�/�/�/*?!? 3?`?W?i?�?�?�?�? �?�?�?�?&OO/O\O SOeOO�O�O�O�O�O �O�O"__+_X_O_a_ {_�_�_�_�_�_�_�_ oo'oToKo]owo�o �o�o�o�o�o�o #PGYs}�� �������L� C�U�o�y�������܏ ӏ��	��H�?�Q� k�u�������؟ϟ� ���D�;�M�g�q� ������ԯ˯ݯ
�� �@�7�I�c�m����� ��пǿٿ����<� 3�E�_�iϖύϟ��� ��������8�/�A� [�eߒ߉ߛ��߿��� �����4�+�=�W�a� ������������� �0�'�9�S�]����� ��������������, #5OY�}�� �����(1 KU�y���� ���$//-/G/Q/ ~/u/�/�/�/�/�/�/ �/ ??)?C?M?z?q? �?�?�?�?�?�?�?O O%O?OIOvOmOO�O �O�O�O�O�O__!_ ;_E_r_i_{_�_�_�_ �_�_�_ooo7oAo noeowo�o�o�o�o�o �o3=ja s������� ��/�9�f�]�o��� ����ҏɏۏ���� +�5�b�Y�k������� Οşן����'�1� ^�U�g�������ʯ�� ӯ ���	�#�-�Z�Q� c�������ƿ��Ͽ�� ���)�V�M�_ό� �ϕ��Ϲ�������� �%�R�I�[߈�ߑ� �ߵ����������!� N�E�W��{���� ����������J�A� S���w����������� ����F=O| s������� B9Kxo� ������// >/5/G/t/k/}/�/�/ �/�/�/�/??:?1? C?p?g?y?�?�?�?�? �?�?�?	O6O-O?OlO cOuO�O�O�O�O�O�O �O_2_)_;_h___q_ �_�_�_�_�_�_�_o .o%o7odo[omo�o�o �o�o�o�o�o�o*! 3`Wi���� ����&��/�\� S�e�������ȏ��я ���"��+�X�O�a� ������ğ��͟�� ��'�T�K�]����� ������ɯ���� #�P�G�Y���}����� ��ſ߿����L� C�Uς�yϋϸϯ��� �����	��H�?�Q� ~�u߇ߴ߽߫����� ���D�;�M�z�q� ���������
�� �@�7�I�v�m���� ����������< 3Eri{��� ���8/A new����� ��/4/+/=/j/a/ s/�/�/�/�/�/�/�/ ?0?'?9?f?]?o?�?|�?�=  �8 �?�?�?OO/OAOSO eOwO�O�O�O�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o �o�o�o�o�o�o# 5GYk}��� ������1�C� U�g�y���������ӏ ���	��-�?�Q�c� u���������ϟ�� ��)�;�M�_�q��� ������˯ݯ��� %�7�I�[�m������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� ��������/�A�S� e�w߉ߛ߭߿����� ����+�=�O�a�s� ������������ �'�9�K�]�o����� ������������# 5GYk}��� ����1C Ugy����� ��	//-/?/Q/c/ u/�/�/�/�/�/�/�/ ??)?;?M?_?q?�? �?�?�?�?�?�?OO %O7OIO[OmOO�O�O �O�O�O�O�O_!_3_ E_W_i_{_�_�_�_�_ �_�_�_oo/oAoSo eowo�o�o�o�o�o�o �o+=Oas �������� �'�9�K�]�o����� ����ɏۏ����#� 5�G�Y�k�}������� şן�����1�C� U�g�y���������ӯ ���	��-�?�Q�c��u���������  ����ٿ���� !�3�E�W�i�{ύϟ� ������������/� A�S�e�w߉ߛ߭߿� ��������+�=�O� a�s��������� ����'�9�K�]�o� ���������������� #5GYk}� ������ 1CUgy��� ����	//-/?/ Q/c/u/�/�/�/�/�/ �/�/??)?;?M?_? q?�?�?�?�?�?�?�? OO%O7OIO[OmOO �O�O�O�O�O�O�O_ !_3_E_W_i_{_�_�_ �_�_�_�_�_oo/o AoSoeowo�o�o�o�o �o�o�o+=O as������ ���'�9�K�]�o� ��������ɏۏ��� �#�5�G�Y�k�}��� ����şן����� 1�C�U�g�y������� ��ӯ���	��-�?� Q�c�u���������Ͽ ����)�;�M�_� qσϕϧϹ������� ��%�7�I�[�m�� �ߣߵ���������� !�3�E�W�i�{��� ������������/� A�S�e�w��������� ������+=O as������ �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?y?�?�?�? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O �O�O__)_;_M___ q_�_�_�_�_�_�_�_ oo%o7oIo[omoo �o�o�o�o�o�o�o !3EWi{�� �������/� A�S�e�w��������� я�����+�=�O� a�s���������͟ߟ ���'�9�K�]�o� ��������ɯۯ��� �#�5�G�Y�k�}���(����ñǰ��ݿ ���%�7�I�[�m� ϑϣϵ��������� �!�3�E�W�i�{ߍ� �߱����������� /�A�S�e�w���� ����������+�=� O�a�s����������� ����'9K] o������� �#5GYk} �������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ������������ /ASew��� ����+= Oas����� ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?5?G?Y?k?}?��?�?�?�9�$FE�AT_DEMOIoN  �4��0���0�4INDE�X�;�1��0IL�ECOMP k����+A��2�5!@SETUPo2 l+E5B?�  N `AC�_AP2BCK �1m+I  �)�8�O�K%�O�O�0.@�O�O�5�O_�O B_�OO_x__�_+_�_ �_a_�_�_o,o�_Po �_to�oo�o9o�o]o �o�o(�oL^�o ���G�k � ��6��Z��g��� ���C�؏�y���� 2�D�ӏh�������-� Q��u�����@� ϟd�v����)���Я _������*���N�ݯ r�����7�̿[�� ϑ�&ϵ�J�\�뿀� Ϥ϶�E���i��ύ� �4���X���|ߎ�� ��A�����w���0� B���f��ߊ�����t:In@PrO 2�@*.VR����*�:�|�@�d�N����PCl����F'R6:����P���t�T	@	��E��0��kM�*.F���~�	���8X�|STM�"���M�q|H>�3�Oa�}
GIF /*/5/p��z/}
JPG�/��/5�/W/i/�/u�JS?1?��#?�/�%
JavaSc�ript]?�/CS�N?�?4�?_? %�Cascadin�g Style ?Sheets�?S��
ARGNAME�.DTOs�8\@$O�?D1TDeOOT@�DISP*[Oq��PD�OiO{A�A�O�O
�TPEINS.X3ML_@O:\,_�O�LACustom Toolbarm_��IPASSWOR�D�Oq�FRS:�\�_o_�@Pass�word Config�_L�:o�_3o po��o#o�o�oYo�o }o$�oH�ol�o �1�U���  ��D�V��z�	��� ��?�ԏc�������.� ��R��K������;� П�q����*�<�˟ `���%���I�ޯ m�ׯ���8�ǯ\�n� ����!���ȿW��{� ϟ���F�տj���c� ��/���S����ω�� ��B�T���x�ߜ�+� =���a��߅���,�� P���t����9��� ��o����(�����^� ����{���G���k�  ��6��Zl�� ��CU�y �D�h��� -�Q���/� @/��v//�/)/�/ �/_/�/�/?*?�/N? �/r?�??�?7?�?[? m?O�?&O�?O\O�? �OO�O�OEO�OiO�O _�O4_�OX_�O�O�_ _�_A_�_�_w_o�_ 0oBo�_fo�_�o�o+o �oOo�oso�o�o> �o7t�'�� ]���(��L���p��������$F�ILE_DGBCK 1m������� �< �)
SUMMARY.DG���\�MD:�$��h�Diag S?ummary%�2��
CONSLOG�����h���7�C�onsole l�og��1�	TPA'CCN���%�(��3�TP Acc?ountinʟ2��FR6:IPKDMP.ZIP\��`�
t���4�D�Exception���b��MEMCHECCK����4����Memory D�ata5���(i{�)�RIPE��p����C�%{�� Packet 9Lɟk��9��{�STAT������<�� %вSt�atus=��	F�TP���#Ϙ�?����mment T�BD��i���)�ETHERNE�ϙ���D�7�E�thernٰ��figuraЯ8���?DCSVRF�ϛ�����M��� ve�rify all���l��|��DIFF�ߤ߶�K�ʳ��diffM����CHG01B�)�;����O�c���o���P��2����T�_������3J�1�C���� j�����VT�RNDIAG.LAS����\G�O Opel�۱ <��nostici���$�)VDEV DAT]:L^�P�VisDe�vice��IM�G ����bɳ��Imag��UP� ES�=�FRS:\���8�Updates� List�2��PFLEXEVEAN:�ASl/O�/! UIF Ev���ܿm����)
P�SRBWLD.C	M�/\���/����PS_ROBOW�EL��0�X GR�APHICS4D�b/K/]/o/%4�D Graphics File^��n��8v�GIG�~��?^?�?B�Gi�gE��/m��`v�SM��RO�?vOA��?A/Email���a"O0E7� hAHADOWrOWOiO�O�E�Shadow? Chang�?j�� ���BRCME�RR�O�O�O�_E��GPCFG Err�or� t�@%_ ���8��CMSGLIBz_a_s_oB��UX�	 �0	o�P�$)�PZDCObo�_܆oA�ZD@ad�(o�\�l�BNOT�I��eowoC�N?otificmҵo�j��}�v�PMIOQo�o�o�FWqOnb��7�RtUI[0m��xUI��7)��l��[���+0Ԁ��Ï*6���� ����8�J�ُn��� ��!�3�ȟW������ "���F�՟?�|���� /�į֯e�������� ��T��x������=� ҿa�˿ϗ�,ϻ�P� b���Ϫ�9�K��� o��ߥ�:���^��� Wߔ�#߸�G�����}� ��6�����l��ߐ� ��1���U���y��� � ��D���h�z�	���-� ��Q�c�����.�� R��vo�;� _��*�N� ����I�m /��8/�\/��/ �/!/�/E/�/i/{/? �/4?F?�/j?�/�?? �?�?S?�?w?OO�? BO�?fO�?O�O+O�O �OaO�O�O_�O_P_ �Ot__�_�_9_�_]_ �_�_�_(o�_Lo^o�_ �oo�o5o�o�oko  �o$6�oZ�o~��ox�$FIL�E_FRSPRT�  ���p�����xM�DONLY 1m��usp 
 ��)MD:_VD�AEXTP.ZZ�Z�qH�W�6�%NO Back file "�9����N��8� ͏�ڏ�H'���K� ]�쏁������F�۟ j������5�ğY�� f������B�ׯ�x� ���1�C�үg����� ��,���P��t��� ��?�οc�u�ϙ�(� ����^��ς��)��t?VISBCK ��q>�*.VD*�t߾��FR:\C�I�ON\DATA\�_�����Vis?ion VDu���~��*.CAM���� %	���ӕߧ��GigE Ca�mera Definit��$��t� �Ϙ��ϑ���]���� �(���L���p���� ��5�����k� ��$ ��Z��~�� C�g��2� Vh���?� �u
/�/@/�d/�.�LUI_CON�FIG n�u�V�s+ $ Q#�{�u�/�/�/ ?0?$?29� |xZ/\? n?�?�?�?�<J?�?�? �?OO�?0OUOgOyO �O�O4O�O�O�O�O	_ _�O?_Q_c_u_�_�_ 0_�_�_�_�_oo�_ ;oMo_oqo�o�o,o�o �o�o�o�o7I [m�(��� ����3�E�W�i� {������ÏՏ��� ���/�A�S�e�w�� ������џ������ +�=�O�a�s�
����� ��ͯ߯񯈯�'�9� K�]�o��������ɿ ۿ���#�5�G�Y� k�Ϗϡϳ�����n� ����1�C�U���y� �ߝ߯�����j���	� �-�?�Q���u��� �����f�����)� ;�M���q��������� ��b���%7I ��m����^ ��!3�Di {���H��� ////�S/e/w/�/ �/�/D/�/�/�/?? +?�/O?a?s?�?�?�? @?�?�?�?OO'O�? KO]OoO�O�O�O8O�O��O�O�O_#_�H � x/_<S�$F�LUI_DATA o���lQ��A^TR�ESULT 2p�lU�P �T��/wizar�d/guided�/steps/ExpertK_�_�_ �_oo&o8oJo\ono��o�j�Cont�inue wit�h G�Pance �o�o�o�o�o#5`GYk}� =R�->QlU�y0a��@��lQ��_ps��+�=�O�a� s���������͏ߏ�` �O��*�<�N�`�r� ��������̟ޟ����"��|�vrip �P�h�z�������¯ ԯ���
��.��R� d�v���������п⿀����*�<���� ��|��v��PTi�meUS/DST D���������&�8��J�\�n߀ߗgEnabl�o�������� ��� �2�D�V�h�z�
��=R�������Ϭ�24���.�@� R�d�v����������� �ߡ�*<N` r�������������#�w�_�QRegion�p�� ����� //$/��kAmerica\�^/p/�/�/�/�/ �/�/�/ ??$?��A�y�n?�?B�Sditor5?�?�?�? �?OO0OBOTOfOxO��kYular  �?�O�O�O�O�O__�1_C_U_g_y_8?� ��� �?d?�_�?�?/accesM/o)o ;oMo_oqo�o�o�o�o��o:�Conne�ct to Network�o# 5GYk}�����B8��_�_�(���!�_�0Introduct\o��� ������ɏۏ���� #�>�G�Y�k�}����� ��şן�����1� N��N�x��_�6updat����ѯ �����+�=�O�a��s�2�Not r�ight now ����ƿؿ���� ��2�D�V�h�z�=<� N?\�����@���	�� -�?�Q�c�u߇ߙ߫� ����:�����)�;� M�_�q�������"�	���Ϭ���� ��C�U�g�y������� ��������	��? Qcu����� ��)����� n0������� //%/7/I/[/m/, ~/�/�/�/�/�/�/? !?3?E?W?i?{?:�? ^�?��?�?OO/O AOSOeOwO�O�O�O�O �O�?�O__+_=_O_ a_s_�_�_�_�_�_�? �_�?o�?9oKo]ooo �o�o�o�o�o�o�o�o #�OGYk}� �������� �_@�od�&o(����� ��ӏ���	��-�?� Q�c�u�4������ϟ ����)�;�M�_� q�0���T���ȯ��� ��%�7�I�[�m�� ������ǿ������ !�3�E�W�i�{ύϟ� ���ς�̯�����ܯ A�S�e�w߉ߛ߭߿� ��������ؿ=�O� a�s��������� ���������B�l� .ߓ������������� #5GYk*� ������ 1CUg&�8�J�\� �����	//-/?/ Q/c/u/�/�/�/�/| �/�/??)?;?M?_? q?�?�?�?�?�?�� �O�7OIO[OmOO �O�O�O�O�O�O�O_ �/3_E_W_i_{_�_�_ �_�_�_�_�_oo�? �? Obo$O�o�o�o�o �o�o�o+=O a _r����� ���'�9�K�]�o� .o��Ro��voۏ��� �#�5�G�Y�k�}��� ����ş֏����� 1�C�U�g�y������� ����⯤��ȏ-�?� Q�c�u���������Ͽ ����֟;�M�_� qσϕϧϹ������� ��ү4���X��� �ߣߵ���������� !�3�E�W�i�(ύ�� ������������/� A�S�e�$߆�Hߪ��� ������+=O as����z�� �'9K]o ����v������ /��5/G/Y/k/}/�/ �/�/�/�/�/�/?� 1?C?U?g?y?�?�?�? �?�?�?�?	O�/� 6O`O"/�O�O�O�O�O �O�O__)_;_M___ ?�_�_�_�_�_�_�_ oo%o7oIo[oO,O >OPO�otO�o�o�o !3EWi{�� �p_�����/� A�S�e�w��������� ~o�o�o��o+�=�O� a�s���������͟ߟ ���'�9�K�]�o� ��������ɯۯ��� �Џ��V��}��� ����ſ׿����� 1�C�U��fϋϝϯ� ��������	��-�?� Q�c�"���F���j��� ������)�;�M�_� q����������� ��%�7�I�[�m�� ������t��������� !3EWi{�� �������/ ASew���� ���/��(/��L/ /�/�/�/�/�/�/ �/??'?9?K?]? �?�?�?�?�?�?�?�? O#O5OGOYO/zO</ �O�Ot?�O�O�O__ 1_C_U_g_y_�_�_�_ n?�_�_�_	oo-o?o Qocouo�o�o�ojO�O �O�o�O);M_ q������� ��_%�7�I�[�m�� ������Ǐُ����o �o*�T�{����� ��ß՟�����/� A�S��w��������� ѯ�����+�=�O� � �2�D���h�Ϳ߿ ���'�9�K�]�o� �ϓϥ�d��������� �#�5�G�Y�k�}ߏ� �߳�r������ߺ�� 1�C�U�g�y���� ����������-�?� Q�c�u����������� ����������J� q������� %7I�Z �������/ !/3/E/W/x/:�/ ^�/�/�/�/??/? A?S?e?w?�?�?�?�/ �?�?�?OO+O=OOO aOsO�O�O�Oh/�O�/ �O�/_'_9_K_]_o_ �_�_�_�_�_�_�_�_ �?#o5oGoYoko}o�o �o�o�o�o�o�o�O �O@_y��� ����	��-�?� Q�ou���������Ϗ ����)�;�M� n�0����h�˟ݟ� ��%�7�I�[�m�� ����b�ǯٯ���� !�3�E�W�i�{����� ^�����̿�����/� A�S�e�wωϛϭϿ� �����ϴ��+�=�O� a�s߅ߗߩ߻����� �߰���Կ�H�
�o� ������������� �#�5�G��k�}��� ������������ 1C��&�8�\� ����	-? Qcu��X��� ��//)/;/M/_/ q/�/�/�/fx��/ �?%?7?I?[?m?? �?�?�?�?�?�?�O !O3OEOWOiO{O�O�O �O�O�O�O�O�/�/�/ >_ ?e_w_�_�_�_�_ �_�_�_oo+o=o�? Noso�o�o�o�o�o�o �o'9K
_l ._�R_����� �#�5�G�Y�k�}��� ���ŏ׏����� 1�C�U�g�y�����\ ���⟤	��-�?� Q�c�u���������ϯ �󯲏�)�;�M�_� q���������˿ݿ� ���ҟ4�����m�� �ϣϵ���������� !�3�E��i�{ߍߟ� ������������/� A� �b�$φ��\߿� ��������+�=�O� a�s�����V߻����� ��'9K]o ��R��v����� #5GYk}� �������// 1/C/U/g/y/�/�/�/ �/�/�/���?<? �c?u?�?�?�?�?�? �?�?OO)O;O�_O qO�O�O�O�O�O�O�O __%_7_�/??,? �_P?�_�_�_�_�_o !o3oEoWoio{o�oLO �o�o�o�o�o/ ASew��Z_l_ ~_��_��+�=�O� a�s���������͏ߏ �o��'�9�K�]�o� ��������ɟ۟ퟬ ��2��Y�k�}��� ����ůׯ����� 1���B�g�y������� ��ӿ���	��-�?� ��`�"���F��Ͻ��� ������)�;�M�_� q߃ߕߦϹ������� ��%�7�I�[�m�� ��Pϲ�t������� !�3�E�W�i�{����� ����������/ ASew���� ������(��� as������ �//'/9/��]/o/ �/�/�/�/�/�/�/�/ ?#?5?�V?z?�? P/�?�?�?�?�?OO 1OCOUOgOyO�OJ/�O �O�O�O�O	__-_?_ Q_c_u_�_F?�?j?�_ �_�?oo)o;oMo_o qo�o�o�o�o�o�o�O %7I[m ������_�_�_ �0��_W�i�{����� ��ÏՏ�����/� �oS�e�w��������� џ�����+��� � ���D�����ͯ߯ ���'�9�K�]�o� ��@�����ɿۿ��� �#�5�G�Y�k�}Ϗ� N�`�r��ϖ����� 1�C�U�g�yߋߝ߯� ���ߒ���	��-�?� Q�c�u������� ��ϲ���&���M�_� q��������������� %��6[m ������� !3��T�x:�� �����//// A/S/e/w/�/��/�/ �/�/�/??+?=?O? a?s?�?D�?h�?� �?OO'O9OKO]OoO �O�O�O�O�O�O�/�O _#_5_G_Y_k_}_�_ �_�_�_�_�?�_�?o �?�_Uogoyo�o�o�o �o�o�o�o	-�O Qcu����� ����)��_J�o n���D����ˏݏ� ��%�7�I�[�m�� >����ǟٟ���� !�3�E�W�i�{�:��� ^���ү������/� A�S�e�w��������� ѿ������+�=�O� a�sυϗϩϻ��ό� ֯����$��K�]�o� �ߓߥ߷��������� �#��G�Y�k�}�� ������������� ������v�8ߝ��� ��������	-? Qcu4���� ��);M_ q�B�T�f����� //%/7/I/[/m// �/�/�/�/��/�/? !?3?E?W?i?{?�?�? �?�?�?���O� AOSOeOwO�O�O�O�O �O�O�O__�/*_O_ a_s_�_�_�_�_�_�_ �_oo'o�?Ho
Olo .O�o�o�o�o�o�o�o #5GYk}�o �������� 1�C�U�g�y�8o��\o ���o���	��-�?� Q�c�u���������ϟ ����)�;�M�_� q���������˯��� ���ҏԯI�[�m�� ������ǿٿ���� !���E�W�i�{ύϟ� ������������ܯ >� �b�t�8ϛ߭߿� ��������+�=�O� a�s�2ϗ������� ����'�9�K�]�o� .�x�Rߜ��������� #5GYk}� ������� 1CUgy��� ��������/��?/ Q/c/u/�/�/�/�/�/ �/�/??�;?M?_? q?�?�?�?�?�?�?�? OO���/jO,/ �O�O�O�O�O�O�O_ !_3_E_W_i_(?�_�_ �_�_�_�_�_oo/o AoSoeowo6OHOZO�o ~O�o�o+=O as����z_� ���'�9�K�]�o� ��������ɏ�o�o�o ��o5�G�Y�k�}��� ����şן����� �C�U�g�y������� ��ӯ���	��ڏ<� ��`�"���������Ͽ ����)�;�M�_� qς��ϧϹ������� ��%�7�I�[�m�,� ��P���t�������� !�3�E�W�i�{��� �����������/� A�S�e�w��������� ~���������=O as������ ���9K]o �������� /��2/��V/h/,�/ �/�/�/�/�/�/?? 1?C?U?g?&�?�?�? �?�?�?�?	OO-O?O QOcO"/l/F/�O�O|/ �O�O__)_;_M___ q_�_�_�_�_x?�_�_ oo%o7oIo[omoo �o�o�otO�O�O�o �O3EWi{�� �������_/� A�S�e�w��������� я�����o�o�o�o ^� ��������͟ߟ ���'�9�K�]�� ��������ɯۯ��� �#�5�G�Y�k�*�<� N���r�׿����� 1�C�U�g�yϋϝϯ� n�������	��-�?� Q�c�u߇ߙ߽߫�|� �����Ŀ)�;�M�_� q����������� ����7�I�[�m�� �������������� ��0��T�{�� �����/ ASev���� ���//+/=/O/ a/ �/D�/h�/�/ �/??'?9?K?]?o? �?�?�?�?v�?�?�? O#O5OGOYOkO}O�O �O�Or/�O�/�O�/�O 1_C_U_g_y_�_�_�_ �_�_�_�_	o�?-o?o Qocouo�o�o�o�o�o �o�o�O&�OJ\  o������� ��%�7�I�[�o� ������Ǐُ���� !�3�E�W�`:�� ��p՟�����/� A�S�e�w�������l� ѯ�����+�=�O� a�s�������h����� ֿ �'�9�K�]�o� �ϓϥϷ��������� ��#�5�G�Y�k�}ߏ� �߳��������ߺ�̿ ޿�R��y���� ��������	��-�?� Q��u����������� ����);M_ �0�B�f���� %7I[m ��b�����/ !/3/E/W/i/{/�/�/ �/p���/�?/? A?S?e?w?�?�?�?�? �?�?�?�O+O=OOO aOsO�O�O�O�O�O�O �O_�/$_�/H_
?o_ �_�_�_�_�_�_�_�_ o#o5oGoYoj_}o�o �o�o�o�o�o�o 1CU_v8_�\_ ����	��-�?� Q�c�u�������joϏ ����)�;�M�_� q�������fȟ�� ���%�7�I�[�m�� ������ǯٯ����� !�3�E�W�i�{����� ��ÿտ������ܟ >�P��wωϛϭϿ� ��������+�=�O� �s߅ߗߩ߻����� ����'�9�K�
�T� .�x��d��������� �#�5�G�Y�k�}��� ��`��������� 1CUgy��\� �������-? Qcu����� ����/)/;/M/_/ q/�/�/�/�/�/�/�/ ����F?m?? �?�?�?�?�?�?�?O !O3OEO/iO{O�O�O �O�O�O�O�O__/_ A_S_?$?6?�_Z?�_ �_�_�_oo+o=oOo aoso�o�oVO�o�o�o �o'9K]o ���d_v_�_��_ �#�5�G�Y�k�}��� ����ŏ׏鏨o��� 1�C�U�g�y������� ��ӟ������<� �c�u���������ϯ ����)�;�M�^� q���������˿ݿ� ��%�7�I��j�,� ��P������������ !�3�E�W�i�{ߍߟ� ^�����������/� A�S�e�w���Zϼ� ~���Ϥ��+�=�O� a�s������������� ����'9K]o ��������� ��2Dk}� ������// 1/C/g/y/�/�/�/ �/�/�/�/	??-??? �H"l?�?X�?�? �?�?OO)O;OMO_O qO�O�OT/�O�O�O�O __%_7_I_[_m__ �_P?�?t?�_�_�?o !o3oEoWoio{o�o�o �o�o�o�o�O/ ASew���� ���_�_�_�_:��_ a�s���������͏ߏ ���'�9��o]�o� ��������ɟ۟��� �#�5�G���*��� N���ůׯ����� 1�C�U�g�y���J��� ��ӿ���	��-�?� Q�c�uχϙ�X�j�|� �Ϡ���)�;�M�_� q߃ߕߧ߹����ߜ� ���%�7�I�[�m�� ������������ ��0���W�i�{����� ����������/ AR�ew���� ���+=�� ^ ��D����� �//'/9/K/]/o/ �/�/R�/�/�/�/�/ ?#?5?G?Y?k?}?�? N�?r�?��?OO 1OCOUOgOyO�O�O�O �O�O�O�/	__-_?_ Q_c_u_�_�_�_�_�_ �_�?o�?&o8o�O_o qo�o�o�o�o�o�o�o %7�O[m �������� !�3��_<oo`���Lo ��ÏՏ�����/� A�S�e�w���H���� џ�����+�=�O� a�s���D���h���ܯ ����'�9�K�]�o� ��������ɿۿ���� �#�5�G�Y�k�}Ϗ� �ϳ����ϖ�����̯ .��U�g�yߋߝ߯� ��������	��-�� Q�c�u������� ������)�;�����߀����$FMR�2_GRP 1q���� ��C4  B�.C�	 C�����^��E�� ���<����P]��P�W��Pm4�M��D$L��?� @<���:N��:�o:I���9-�tA��  ��BH��C���NC�  C����h�<��������@UUU�UU�I��>��$�<�6=�¹�=f'�=�m�=���;:�;:,��:���: �:�7�:��� (�L���/��//B��_CFG {r��T :/�{/�/�/A+NO ���F268�925   @,R�M_CHKTYP  ��C�������ROM� _MI9N� C���"0��X��SSBQ#s��� ���O?C�F3o?�?G%T�P_DEF_OW�  C���7I�RCOM� �?�$�GENOVRD_�DO6M��=TH�R6 d�5d�4_�ENB�? �0RWAVC��t87C0� ���@ E�#	�E
��F�� FZ\�FC��?%/�OC���#0�E�O���B�:AOU��z����!���2��<0R,_�O$_F_t_C�C�� ��_U0�_�]@�]B���Rp��Y�?;@SMT���{HI��E0�T�$HoOSTCQ"1|��nD0�M� 	ohMokooC��o@�e�o�o�o" ?��oSew��o��@pr01 ymous�����&� no�o�oo���o B��ɏۏ�4�#��5�G�Y�|���wilder ����� ̟ޟ�7�I�[�8�o� \�����������}�s������"�E�F� e	anon�q��� ������ ��$�6�8� %�l�I�[�m�ϑ�د �����������V�3� E�W�i�{�¿����� ���.����/�A�S� ��w�������� *���+�=�O��ߨ� ������������ 'n�K]o�� ��������# j�|���k���>� ���0//1/C/ U/x���/�/�/�/ �/,>Pbd/Q?� u?�?�?�?�?/�?�? OO)OL?�/�/qO�O�O�O�OMeENT �1}�K P!�? omput���O�g`�@72.22.19.4 _ b�@=_O_Ui_,_�_ �_b_�_�_�_�_o�_ /o�_oeo(o�oLo�o po�o�o�o�o+�o Os6lZ�� �����9��]� o�2���V���z�ۏ�� ��ԏ5���Y��}��@���d�v�ן !?QUICC0ٟ���!19P68.?10.201 �閼&��!1V136P��2y�U�ǟ�ȯ!ROUTERɯ��!�B���?PCJOG����f���0��CAMPRTi�E�� ���w�RT⯔����� !Softw�are Oper�ator Pan�el�V�W��DNA�ME !�J!�ROBO��_�S_�CFG 1|�I� �Au�to-start{ed4FTP?��2?4O�h??�Q� c�u߇��?�߽����� ��ߘ�)�;�M�_�q� �.���������#��� �$�6�H��l�~��� ������Y����� �2D�'
ROS_�I Tag�	SM?�����&9�� ����7I[ m�$����,�/*�Xg��t �c/���/�/�/�/ �/�??)?;?M?p/��/�?�?�?�?�?.����wilder-�@/R//Of?�/QO wO�O�O�Ot?�O�O�O __<O�OO_a_s_�_�_.��>��OO�_ 2_TOoCoUogoyo@_ �o�o�o�o�oo�o -?Qc.��� 	�x�X+b�_�o� ����+�=�O�s� ���������`��� �'�9���口��� ɏ���ڟ����׏ 4�F�X�j�|���!����į֯������_ERR ~x��&��PDUSIZ  ���^Ő�=�>~V�WRD ?���,a�  �abc t����gues����п����k�SCDMNG�RP 2��@�����������K5� 	P0�2.00 8�� o  8��i���  
�q�� � �c� �������
��:����U�����i�}��P`�P�m�	�~}����������0���  e�i��q�8�
+q�����~���!���"�����ՙ��V���s�GY��aׂ��da�sυϗ��_�GROU ��5��7���	�01.�0k��QUPD � (e=���	�T�Y��5�(�TT�P_AUTH 1��5� <!i?Pendan��r������ !K?AREL:*r�{���KC�������VISION �SET��"����V! 9�'�Q���u�c������������
����A�C?TRL �5�P��[
  �?FFF9E3���FRS:DEF�AULT�F�ANUC Web Server�� n 7��D�~���)��,>P$�WR�_CONFIG ;�$� o�&��IDL_CPU_kPC� ��BȎ��� B��v�M�IN�n� >���t�GNR_IO�/�d���;��NPT_SIM_DO��+STAL_S�CRN� ��I�NTPMODNT�OL:'+�RTY�(�&�E�ENB�:'��OLNK 1�5����/�/��/ ??$?6?�"MA�STE��!SL?AVE �5��$�SRAMCACH�ET?f3G�O_CF0\И>�"�3UO,�?~�2CMT_OP� 8�9��3YCL�?�5�� _ASG 1�$�p�
 8?[OmO O�O�O�O�O�O�O�O�_!_3_E_@;.BNU��Pe�9�
�2IP��?�7RTRY_C�N�?�56!&�c��!�b=� �2�0�2�t>���o���P_ME�MBERS 2��$�a� $�Ab���(:g@oRi�RC�A_ACC 2����  U��� g �� )� 6
��-���f�@ �'�~�o�d�x���l�dBUF0���2���= I wu2 "pI u�Яu1I@+t`#t��+t�+t�#t�+sJ�.p]r #sJ2tJ`�[t�ktJtJ�[t�j#sKbtK*tK@�t�ztKBtK��t�tK�ZtL"tL*tL2tL�:tLBtLJtLRtL�ZtMbt(n� � n�Hu� u�Bh#��u2�^j�u1+q��K��u2#q-K�(c�H[�:��e��c��1�1�o  F�K�Fۓ�m�[�GK�G;���[u2T� pG�{u1�U�H� 	��	`H*tH��tHztHBtH�tH�tHZt y21 CUgy��������	���m�"1�dn�9�:P:�I�[�m����𣏵���1	D(xɁˁс^��ُ����s3�(�   2�9�;�9�C�9�K�9�`S�9�[�9�c�  j� q�s�q�D���q���q� \���q���J�=���J� ��J���ʓJ�ӒJ����  ��<���� L�
��\���l�!� a�*�a�2�a�:�a�B� 7�S�7�[�7�c�G�k� G�s�G�{�G�LĊ�G� ��sњ��£��«�s� ���²��º���s� Ƀأ��Ĵ�ؠT����ؠ��
���a�12����4�9�s�s�<�s�U�X���dHIuS
r��� ܠa� 2022-1�2-26�� 
�`�`P_�����߀����/�A�S�U��M ��>����P� + �P %� '��+�H  � *�PF(��-��  ( !X�H   0 mP	 3���������X�0�g�Um�0z��  ;Z�c� ; ���g�� . #   &����8��# )@ �� >�� '3 #�0��"U��<%���������c�7�= ��09-2z��� �����e�U�m�0�l�L������Z�c��<��f�U6�`&�ڪ�P���P,[�J��4�PW��"  8����U�XВ�_  0��#<w;B��� ?��s����~�;�`U5 yꔸP.m�NU�X�d���9�`_��0 2�����.I@��+�LF/X/j/|/�,� �  5 
� 6� Y�!"U0D�&16V�Xй�X�r�@E^X�Bi����,D� /@ �0? -???Q?c?u?XZp��|ߎߠډ��?�?�? OO0OBOTOfOxOf�Jx�L3�Psb���)!^��!Z��6 G \��]��4+mP��__,_>_PP_>�P��P
��j�@M��"��!"��7�A���2��T��1��Q�����G0-V��/�@OY_�_oo&o�&805oX��PU�!8 7n '��Aqo�o�o�o�o�o�#��<�  )s �|�, hЩ0�Q�D_��$��;T����=U�����P5��bZ(��C ������2�BrP��"�X0�PR(!"��)�@E���R>  �R)�|������/��� @!"�/�/�/�/�,�����$cq09  a��P�b�t�����@�?s���?�?���������1�C�U�g�`y������Ox����� ���� �����  �<�(� �T�-��
,�������M����1�C�U�g�y�g_T��=٘�c��ܤ���  �ݘ�# ʽ��8 ���@w ��� ����P ���U ����#�5�G�Y�GoF4	�� �T	��0��0������������߾��� ��#ƪU�Ԥ�ܤ����죣�Ǭć�ܰ���<�B��ҼϹ���������8��<ѿ` ����G�ƨ��c��ܰ�വ��I�@��N����ﳏ�	�<�8м�g�ۏƪ�Ԥ���İ��P���ܰ�ഔ<�D�ʦ��q�������������I_CF�G 2�Ǜ H�
Cycle �TimeB�usy��Idylmin�>uUp	�Read�Dow0,;�A���Count		ONum ������д�1PROG����Ǖѐ��)/softpa�rt/genli�nk?curre�nt=menup�age,1133,ç#5GY4���SDT_ISOL�C  Ǚ��`���J23_DSP_ENB  ��0�INC ���{S�AWp?� � =���<#�y
��:�o�P��./{T/Y/�OB�� C���<�s!G�_GROUP 1푓�R< �� ���/a/�I��/{PQ?9?K?�]??�?�?�?�?���I/k)G_IN_A�UT�P����PO�SRE{/�&KANJI_MASKF�JKARELMO�N �Ǜ�{Ry |?�O�O�O�O�O��SBJ����{T�E|O�KCL_L�0�NUM�4_$KE�YLOGGING��p̐��Q�� LA�NGUAGE �Ǖ�P�DEFAULT �Q6��LD����	YP?pc�PG�R��
<��xhpÀnq�[���'��  /� 
�끛��3�;��
Va(?UT1:\�Ovo �p�o�o�o�o�o�o�o �o(:c�O��5�PN_DISP ��9??>�TOCTOL�p��Dz�����qGB�OOK ��]d`_t�bqbq3�XBl W�i�{���������c=Ӊ��	��Y�!�r�<n�_BU�FF 2�� �c�W�b�2�w ~�6����ٟП�� ��E�<�N�{�r��� ����կ̯ޯ��t� ?DCS ��]" Ќ�����s��������"�IO 2��[C ��޿������ ���*�:�L�^�r� �ϔϦϺ�������� �$�6�J�Z�l�~ߒ�~��ER_ITM�d�?�����!�3�E� W�i�{�������� ������/�A�S��wN��SEV�0���TYP��߻���8��b�ARSTR_ ��SCRN_FL +2�˽��S�S�ew������T�PhP����}NG�NAM�L��R�tU�PS�pGI E��._LOAD�x G %�
%��1_CALIB_�DRIL�~�MAXUALRMOR,?Aۀ��
�4'_PR9?@ �с��B_PNP_D�v�2��	M�DR0771Yuz�"�8063΃@ �#�Yr%/�C�p��_�����o�U#_GRP 2]�#� �r�	�+� Z ;|/6% �� ?�/$?@j?U?? y?�?n?�?�?�?�?�? 	O�?-OOQOcOFO�O rO�O�O�O�O�O_�O )_;____J_�_n_�_ �_�_�_�_oo�_7o "o[oFoo�oto�o�o �o�o�o�o3W iL�x���� ���/�A�$�e�P� ����~������Ώ�����=�(�a��DBGDEF �^%�k!j!l�~�_LDX�DISA���M�EMO_APE� ?�
  >,����"�4�F�X��j��FRQ_CF�G �^'��AM d�@���4 <k$Cd%>/ܯ���"�^+��$*z"�/$� **:-� 4$ �2�˯4&X�j��� ����ͿĿֿ�O�^%�,Ϣ��S�A�v�`�,(Ϫ�4$���ϼ��� ��
�/��S�:�w߉� p߭ߔ��������?ISC 1��	� �l�O��$��e�P��������%�_MS�TR �{���S_CD 1�۝��� 4���X�C�|�g����� ����������	B -Rxc���� ���>)b M�q����� /�(//L/7/p/[/ m/�/�/�/�/�/�/? �/"?H?3?l?W?�?{? �?�?�?�?�?O�?2O OVOAOzOeO�O�O�O �O�O�O�O__@_��MK�����šR_$MLTARM�����}R �FÎ��_�T}�METsPU��3R�����NDSP_ADC�OL�U���^CMNmT�_ �UFN`|o�WFSTLI@o1g�� ���n�S�š�o�d�UPOSC�Fag*nPRPMlo�iST�P1���w 4��#�
/q D�/u?Mw+MOa �������� �E�'�9�{�]�o�������QSING_C�HK  Co$M7ODA���-�{[�}Y�DEV }	��	MC:��>�HSIZE��3P���TASK �%��%$1234?56789 ������TRIG 1��� l}�ʯ�L�0ڟ�L�n�YPY�L����EM_IN�F 1��`�)AT&FV0�E0 ���)�E�0V1&A3&B�1&D2&S0&�C1S0=��)GATZ���ҤH� ����?�ΨAG�o� *���z���ɿ }�� ����ůׯH���lϣ� �Ϣ�U��ρ�������  �ӿ�V�	��-Ϟ� ��c�����߽߳�.� ��R�9�v��;߬�_� q߃ߕ����*�a�;� `���?��������� ���������\n !�����q{��� �4F��j/ AS�w��1/ �B/�S/x/_/�/U^�ONITOR|`G� ?3�   	?EXEC17S�"U2�(3�(4�(5�(T���&7�(8�(97S�"fJ4�"J4�"J4 �"J42J42J4 2J4@,2J482J4D2J32Q8U2]82i82u82�8U2�82�82�82�8U2�83Q83]83�"��R_GRP_S�V 1�l� (����:B����#����?ԡ�c?q�齫G��Ĵ�&�)v�_�D;"\��CION_�DB�����3Q � �3P���E���K�3P�`�� N� �`,3�KO�-ud1E�[_m__�Q�PL_NAME �!}��P�!�R-2000iC�/210L, H�andlingT�ool  *Q�QR�R2cA 1�?�H���Q P\ d�b�_oo +o=oOoaoso�o�o�o �o�o�o�o'9K]o�2�_�� ������*�<�R�f�x������� ��ҏ�����,�>� P�b�t���������Ο �����(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�~� ������ƿؿ���π �2�D�V�h�zωP< U��ϴ����������  �2�D�V�h߅Y��JR �Ϣ�
���߉TP������(�:�L� ^�p��������� �� �����6�H�Z�l� ~���������������  2D�%�z� ������
�.@Rdv��� E@ E5�m��W@  ����Rd��� 
-�,/:'���Z$#�q/�-l/�/� ��(�/�*A�  A=��#�����/�/�?	7�*P�*Q0BH!?��_5�@m?4�@�R�%	`�/�?��?�?�1:�oA �R�?�?Ov�E0*P3B�H0G6$#JQ�� j�P�Pɇ/ �P@嵅��Pv@
<  g�T�E�/�O�/��O�O�O_�O)_�_R�R�S��YL@�2� � �2�lQ @D�  "�Q?��QlQ?^ �Q�^@_f�E;�� �QL�9_  ;��	l�R	 L���X���M@N@�P&�X^,^�X ��R�K����K�3K��1gK���K����K(�.G�}��_�HoRd�=`?�?���?��N@
y�tb�PC���,o� �N����
��ՙ�m`���X�a�4@~3j�9  �p�`�k�ô�`�P�a���k^�� �￑^� �	M�oRr�+s�W�I�O=ogx � �|r_�Yu	�'� � �r�I� �  ��� �PTy:��È�È=�s���u\r@ ��� �pUzrQ*�  L�^rRGH[�Q~9N@0��  '{p���]p@�`?��@/I�@m`@�`���B�[C�`B� ' C4ր�`B�P܂���^ ��CR~"i��	+n� �\ƈ@00�3F4A`� 'I�aX�^Dz_ {�_������՟�v�q�
�` �� �	���q����  �^: 7PC�? ?�ffK/6�H�ڟ �0}���]q8^ �����Q(qȤWw(^ ��q�	���%ax�S�TJ�?333i��]p;���;`H��;S��;�d��;��Y;��*@ܬ�!o[�?X�RrS�R0@?ff�f?�`?&��YtA�#@���@�|g@Բ��� ?Y�����Xu�U迆W �v��Tg�<�'�`�K� ��oϨϓ��������?X�F@0��>��πb�ٿ����U߶�Q�D�a�P��E"� D�߻�	���-�� Q�<�u�`������ EJ��i���_y�?��� f����������_��� ����>)bM�1A���!I���A\�XS��Ul`����/?Y�ز�c��`DC��P��` C�Ї.�	��	����l����Cl�	C~���B41�B���@eaFDÇ�����F�g�p��� ڻ���=�boD��ק��������Y�BG���[�3��:�.�ki_�Y�������B.������m!�D�K�Q�J���L��I�?HخMFEhYt�L.0�LK�F�L��tH���H�0�FE�����!$aLS5��J�G"H�4
H���F�� ��/�/??=?(?a? L?�?p?�?�?�?�?�? O�?'OO7O]OHO�O lO�O�O�O�O�O�O�O #__G_2_k_V_�_z_ �_�_�_�_�_o�_1o oUo@oRo�ovo�o�o �o�o�o�o-Q <u`�����p����Gϭ��%� C�a�M� �ĉ����P�i}�q�����=���� 1�����5��ُ^�y	�� �VwO_������� ��0'�������3&,8����̒Z�؟�����3Xl���@�x�?��3�g�0�0�p�@^����������PP�	P����f��0I�4�m�X�s�z�������ÿҿ�?  I쿮�7� "�[�F��&���Ϡ�����}�������.����1��� ��X�ߠ�����߲�����  2� Eb�E52�mY�B�� �֕ C�~�  @c�^� *�}����p�����#	��
�����#�5��T?�R������ � w����
 B������� ������#5GY`k}�����ԛ����$MR�_CABLE 2��Ԩ Ț�T �@bb?P*�b��Ç����B�C��O4>��B���ߢpH����J�H̼�B�㘤J���,/  ��2�(2�+��  N�/HB�[����g��I�?C��\���CU<``2���^���Bǭ}k���0?h�C����� �.�� ب��/� / /2/�/�/h/�/�/ �/?�/�/�/�/
?? .?�?�?d?�?.�vJ��ۡ B���7��v�;O"O��7�1�
 ����@���� �������@������Y@� ������`�� ��]@U�a@�e@�Y@�m@����`�*�C �D�D�OM� ��	����� �� ?��%% 2345?678901�O�E! �O_�AJ��J�M�ӑJ�
�G�=�not sen�t�JJ�ӐWܥ�TESTFEC�SALGR  e�g��M�d�Ts�1Q
�T�� ��\�J���_�_�_�_ 9U�D1:\main�tenancesG.xmk>o����J��DEFA�ULT���GRP� 2��J  ��PP�p����  ��%!1st c�leaning �of cont.� vYPilati_on 56�R��c!��a�op�+Ǡ���"4FXOn�c%��amech�`cal checki
����sU�q�p�����mv~�aroller���{�����Џ��1�qBasi�c quarte�rlyV�i�{�z,���h�z�������wy�M��J�"8��J� ��p�_�4�F�X�j���˒CM�����ʯ	v#���
��.��}�rGrease� bal0ar b�ush=�����p��篼�ο��A�rCVӐge�r.^�t��y�  3v`D�*�L�S�p�	���ϒ�P�϶���q�gY�,��J�f��-J���p�o�D�V�h�z���q�cabl��J���ӳ���� �
3���,�>�P�@��c)�����|�����������qO?verhauٟ���R� x`\�c�V������������`$�� �4	bi ��Ugy����� "4�-?Q c������� �//f(/M/�P/ ��/�/�/�/�/,/? ?b/7?�/[?m??�? �?�/�??(?�?L?!O 3OEOWOiO�?�O�?�? �OO�O�O__/_~O S_�O�O�_�O�_�_�_ �_�_D_oh_z_Oo�_ so�o�o�o�o
o�o.o @oRodo9K]o� �o��o��� #�5�G��k���� ��ŏ׏���J��1� ��4���y��������� ����F��j�?�Q� c�u���֟������ 0���)�;�M���q� ��ү����˿ݿ�� �b�7φ���mϼ��� �ϵ�����(���L�^� 3߂�W�i�{ߍߟ��� ���$�6�H��/�A� S�e�߉������߽�`������+� /���	 X<�1?��33?�I�>��= �.�&�<2��p��>#�
n�>��OA��B�f�f?L�[-�B �  =�+?��z�?t��=d��f>�a���o<C�;>��q��>��E�n�?'�A7�Y<���͎�����9X?���>�bN>��7>ޯ�z��p�=���m;�D�?��s�n�@@1'A�������q�n���y�#?�?A�>j~�������ѷ>`'R�=�$<�!�-�A!�A��Ũ��-�M��bM��>��y^���P=o>��=�e�z
��XD�B����>��?Co���@  ��P�=	7L>{�6�>�Q���mK �HYk}��C� ����//*/�~N/   ����?+p� K��Q�K��EK����K�OK���eK���K��L%K���K���K���K��%K�Z�K����K�EK��W�K��K�� eK�T�K���%K���r!����� �����`��
 ����@���� � �����@������� �� �����`�� ���� �� ��2�025/12 *>$9 F�@ f/x/ �/�/�/�/�/�/�/? 7��2?D?V?h?z?�? �?�?�?�?�?�?
OO .O@OROdOvO�O�O�O�O�C���ID5U�Q/�_�_�_p�7Q�`�_o0oBop�*5 �_�O�O�O__0_B_�T_f_x_�_�XK p���$MR_HIST� 2���bp� �
 \v�$ 23�45678901PrztHoVbq9o� ����m�+�=�O� ��������`�r��� ����'�ޏK�]�� ��8�����n�۟���� �ȟ5��Y�k�"����F���ů|�鯡�NpS�KCFMAP  ���ep �Ft����ONREL  F��K �EXC/FENBL�
� ��e�FNCl�^�JO�GOVLIML�d�bs���KEYL�z����_PANK��Ӳϲ�RUN������SFSPD�TYP��W��SI�GNL�^�T1MO�T��[��_CE_GRP 1����jrF� ��Ϻ� ����E�����/�A� ��e��uߛ�R߿�v� ���߬��+��O�� s��l��`������ �����9���]�H��PD_THRSH�D  nb@ �w�QZ_EDIT�I��=�TCOM_�CFG 1���o����� 
��_/ARC_i�F���T_MN_MOD�EI���_SP�L%z�UAP_C�PLf{�NOCH�ECK ?� � ��� �'9K]o������5�NO_WAIT_LH����}�ODRDSP�eK�w�OFFSET_CAR��+;&�DISH/9#S_A�@ ARKIǴ�OPEN_FILEg ���� OPTION_IOɿ۱� �M_PRG %��%$$:?^d�!WmO� �(�Ip��:6|d�����'���U0s���U1	 ����U1���� R�G_DSBL  �Zw� ��?8�ORIENTTOK�f��C�*��A 9"�U` IM_D�'���2 V LCT ����N4@Iz��dG_PEXH �j/]DRATH d�w�]D@ UP )�$Ngp����O�O��O�OY�$PAR�AM2�ñ��H��C\W@U�K_]_o_�_�_ �_�_�_�_�_�_o#o 5oGoYoko}o�o�o�o��29_�o�o*@<N`r�/�o �������,� >�P�b�t��������� Ώ�����(�:�L� ^�p���������ʟܟ � ��$�6�H�Z�l� ~�������Ưد��� � �2�D�V�h�z�������¿�<���� � �2�D�V�h�zό� �ϰ��ڰ!�ٿ���@����P��:�L� ^�p߂ߔߦ߸����� �� ��$�6�H��)� ~������������ � �2�D�V�h�z��� [�m���������
 .@Rdv���H������	��!SD� @ R6t���l������0�/~�A�  A�#����//[/Q'e��0��0c!BHi/���%� �/:C  �	`��/�/<?�!:�o�1.?0@?R?d?�B�0{2А �&l���� j������ �@���פ0�0
<  g�4�5��?� O)OOMO8OqO�lT�POU"P�!�_,!��.T�" � �"��A @D� M �A?��C�A?��t�A��C� E;��B��u�O  ;�	l��B	 L���X����0��P&X�^,^X� �BRH����H��cH�DD�H�*sH�_��H<G6G�}�_	�_�T�PBҁ0��0��0�0�Q��AC���x_ ��9  �p�P�k�ùP��@�Q�s4@�_�_ ��[�����Q��=����&��_eB\obb�AwcdG�9�?��_�h  ���bdO�o�e	'� ��  rI� ��  �� ��P�i=���8$6{�b@LRp� Fp�j�Av  L���ǾB�8��nN� �  '�`�t�`-C`B��@4�@�Q��@ ��~[���� � ��CRnY_��	+j^�l�\�� |�{6|14 o9�Q����Dz]OǏYO��֏��!��f�a
��` �� 	�H�qA�A�  Ȇ��:�EsQ�1�@ ?�ff������&� � ɟۛ�a8�������Ata��g( ��-�q9�U�A�qQ,S<,T�s?333�v�`�;���;`H��;S��;�d��;��Y;��*@ܬY�m_�����B��C�Bx0?fff�?�P?&ޠ�dA�#@���@�?|g@Բ����� H�١�F�g�E4��GS� §T����s�����п ����߿�*��N�`� 7τ�oϨ��A�C��Ϭߝ�Da�@��CE"� D�
��U� @�y�dߝ߈��߬��� �����:7�y	��O �ϋ��ϲ�%������� ���!�3���f�Q���hu�����+1A��� 4!��
�������k���?��;B{,f�Y���S�`�]{C��@�` C!Ј�z�U�U T�@�Iܸ���C�l�	C~��B�41�B��@�eaF�^������F�gp���� ڻ��=��bo�]�ק��������Y��BG���[�3��:�Xki_��Y��þ���B.�������m!��]K�Q��J��L���I�Hخ�MFEfX�dL.0��LK�FL���tH���H�0ϺFE�1��$a�LS5�J�G�"H�4
H���F��A/,/ e/P/�/t/�/�/�/�/ �/?�/+??O?:?s? ^?�?�?�?�?�?�?�? O O9O$O6OoOZO�O ~O�O�O�O�O�O_�O 5_ _Y_D_}_h_�_�_ �_�_�_�_�_o
oCo .oSoyodo�o�o�o�o �o�o	�o?*c�N{Gϭkq C�a��� ĉ�8k���~i}q���=�X�}�K�6� [���<%���	4�% ϳVwO��d���<܅l��0'̏ޏ[3&,��
���Z�$�6�����3XlP�b�@��x�?˷3�g�|�|�������Ο(��-P��P6�Q�R�_���k�����������Ư��������0�?  I8�����n������˿r�D����"���� *�4�j�X�z���G�}�g�� ����f���������4�B�  2 EY�[E5^�m���[B�������C�� ��[@��߼�@��������3¿�?�Q�c�u��[?�P��*0�$[[�/�(3[
 ������'�9�K� ]�o��������������Z+�� �����$PARAM�_MENU ?�|�� � DEFP�ULSE��	W�AITTMOUT�?RCVR �SHELL_W�RK.$CUR_oSTYL= ~�OPT�єPTB���CyR_DECSNJ '���� A<N`���������/S�SREL_ID � x����(%US�E_PROG �%#
%/z/)#CC�RV :"��+�'_H�OST !#
!�$�/�*TG��/�#Ĳ/�!�#'?�+_TGIMET:&�% ?GDEBUG8 #�)#GINP_FLgMSKP?9TR�?�7PGA�0 o<�.�;CH�?~8TY+PE ,�// DOmOhOzO�O�O�O�O �O�O�O
__E_@_R_ d_�_�_�_�_�_�_�_ �_oo*o<oeo`oro��o�o�o�o�o�o�5W�ORD ?	#
? 	PRl0���MAI� ��SU�0sTE0���hs	�=rCOL�uhYy}�6LV  }��G�Ȣ%dd1TRA�CECTL 1�v|�- ��7� �S�v 2@��n� �t�2�p�� p� q�2�rDT �Q�|�!��pD� � hN�.���4���4��04�P��4���4�9H�&�S^�1�98�9@� 1�C�U�g�y�������D���9���ം��	⁾�Џ�􏮏@� R�d�v���������П �����*�<�N�`� r���������̯ޯ� "�4����"�4�F�X� j�|�������Ŀֿ� ����0�B�T�f�x� �ϜϮ���������� �,��xߊߜ߮�@�@R�d�����*�N�`��r������� ������&�8�J�\� n��������������� ��"4FXj| ������� 0BTfx�� �����/"/4/ F/X/j/|/�/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?OO,O>OPObOtO�O�On�i,�O�O�O �O__+_=_O_a_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o �o�o�o�o�o�o# 5GYk}��� �����&�8�J� \�n���������ȏڏ ����"�4�F�X�j� |�������ğ֟��� ��0�B�T�f�x���@������ү�OR�j, ��'�9�K�]�o��� ������ɿۿ���� #�5�G�Y�k�}Ϗϡ� ������������1� C�U�g�yߋߝ߯��� ������	��-�?�Q� j�|���������� ����0�B�T�f�x� �������������� ,>Pbt�� ������"a,GYk}� ������// 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O qO�O�N�O�O�O�O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�o�o $6�HZ0f ] W �p^�t_�tՇ�t��t��rg U)�t*�t+�t�tU�t�t�t�tU�t�t�p�F�g�A�r�t�t��t�t�t�t��t	�t
�t�t��t�t�t�t��t�t�t�t*�t�t�t�����z�q �t!�t"��t#�t$�t%�t&J�t'�t(�t�f�Uf$�f,�f4�f��Uf��f��fĄf��f�tf4�f<�f U6�t7�t>�t?�t�@�tA�tB�q� ���	��-�?�Q� c�u���������Ϗ� �����ȯگ� ��*�<�N�`�r�5�Uf<�fD�fL�fT�f\�fd�fl��� '�9�K�]�o������� ��ɿs���������͝UF�tG�tN�tO�tUU�tV�tW�tX�tUY�tZ�t[�t\�q��$PGTRAC�ELEuЅ��A�_�hp����_UP ����������ѬA����_CFG Ȧ����hq	�������A7�C�5�m���C��DEFSP/D ��gq�@����H_CON?FIG �����YD�� d����� gq��PR�5���hp���IN	�T�RL ��1�8lR���PE��ͧ������C���LID
���M�J��LLB 1ϧ�� ���B��B	4��C�$���������E� << fq?��������� A'Iw]�� ������+H��_Vh��������/G�GRP� 1�|��iqCR  �.�hq�B8M�IБ �I״�I�`�Ai�D	6�@������n)~)��E��`L� /��g�.´�#�/�+B� �!�/�/�/�?�/5?hqA� �A�ԚS?�?�>�? <,1�1�?�? �?�?O�?6O!O�?EO@~OAO�O�O�OY z�C�Ohp
�O
_�O_@_ +_d_O_�_s_�_�_�_ �_�_o�_*ooNo��=� )
V7.�10betajE��@�@a?G�@333;!�a�Ci��bf�cDԀ� �ba�cE> �E0� D�` �;!BH��ҡ`< C8����� @��5 �oP�5;!W!�mA�o
q0p�K2��Se<w�  �Do &?@oF6������L�b��-�4�D�e� �u���4�l�~�5�a�p1��CrP� Bq� ɏ���b�`O�}������܄���O�������>�^+���<����;6�V�;E����	t�M���C�ԼB���[�������rW!A*������z3@���������ښ����a������5L�K?NOW_M ��P�|�L�SV է������O������ �ӯ��Я	���v-K�uM#֧� ��b�	0�����	`M��v��V� �����P�@i�ai೵��X�� L�MR#�>�TC9C-�cr��z��K5%�7�-OADB�ANFWD@�J�S�T!1 1���y�47���Ű�P� �ϧϹ��������3� %�7�|�[�m߲ߑߣ� ����������T�3�E�W�v�2��J�����G�<���}�3��������v�4����1�v�5N�`�r���v�A6��������v�7��*v�8GYk�}v�MAa�w$����OVLD  ��m�	/x�PARNUM  �˸1w�SCH�	 �
�L�oãUPDL�%���_CMP_4�� ���p�'m�$ER_wCHK%��m�0V�'&/"+RS �d�N3�_MOaτ(_q/~��_RES_G��ٝ
�b�/<�?�/ +??0?a?T?�?x?�? �?�?�?�?O��#���,�/O�%��.OMO RO�#M�mO�O�O�#�� �O�O�O�#���O
__ �#F *_I_N_�#� i_x�_�_�"V 1ڇ�|v�J��P�\�"THR_INR ����m�d�VMASmS	o ZgMNo�;cMON_QUEUE ۄ�m�J��Pq��N
 UN!N8Kfth�cEND�a�/��iEXE�o�e�B�E<p�o�cOPTI�O�g�+�`PROG�RAM %nj%��`�_r�bTAS�K_I� ~OCFG �no`b�p�DATA7�ݞ{	�e�2����)� ;�M��q����������d�ݏ����~IN+FO7���}�}dΏ k�}�������şן� ����1�C�U�g�y����������ӯ.�:����| �9�q�K_Ƙq��yZ��EN!B� $���D�2M�_��G�q2�$� X�,		X!=��M«���׵ñ$���X!ùù�T�_EDIT ��+�>�tWERFL�h�S�s�RGADJ ���A�  v�?@�0��aZƎa��R��?� ' Bz/��q<ñ�00�%���N��=���2��L�	H�`l���RBpx���Ű��R�*f�/h� **:q�a�s����B�Px���P߀z�������R�Y���DqǼ���4������QBԹPAUUV@(�R��^�p� ���������� �*�x�6���T��F�A�PD������� �����4 �pj|���� ��b^HBT �x����:/� 6/ //,/�/P/�/�/ �/�/?�/?�/�/? ~?(?z?d?^?p?�?�? �?�?�?�?VO ORO<O 6OHO�OlO�O�O�O�O�._�O*___ _J�	���_�p�_�_�T�t$ �_k�_1o�_Uo�go��PREF ��ʄp�p
Z�I�ORITYwƀ>^�MPDSPqLʌ0��gUT�vB�Y�OoDUCT}q��jo�OG�_T�GI��r�rHIB�IT_DOJ�M{TOENT 1��� (!AF_�INE�`��w!�tcI���{!�ud��~!�icm���rXYڝ�����a)�a ~�^�p��`�X� ��|���ŏ���Џ� ��C�*�g�y�`���H����ӟ* s�����0����(�M�>�%��~�/���z��M�����A��,  �`�ïկP���Pş�j�Zj��9�K�]�o�M��E�NHANCE )����A
�di�Ͽ���  ��f�d��o�cT�^�POR_T_NUM�c�`��e^�_CAR�TRE��C�3�S�KSTA�gl{SL�GS�p�C����ó`Unothing׿������������!�3�%{�TEMP �yD�yU� �_a_seiban>o��:o���� �����%��I�4�m� X�j���������� ����E�0�i�T��� x������������� /S>wb�� �����= (:s^���� ���/ /9/$/]/�H/�/l/�/F�{�VE�RSI�`w�  �disabl�e鰼-SAVE ��z	267_0H727�(�/�<?!��>?P?�t? !	�8�b{_�;�?�c�e�?OO+O=OKJ��<s?~O��'_;p �1�C�)0 	�DW�O�OBW^|`URGE��BApe~4�WFPaq�d����fW�p.T�a2�WR�UP_DELAY� �K�0�WR_?HOT %u�b����_?UR_NORMAL�Xr�_�_�WSEMI�_�_6oza_QSKIP�C����Cx�/{o�%����m���et���95�S�������c$ 	Fa�t��?b�C�z�~��D��?j���?��Ģ��8��o�gja�o .@dR��� r�����*�� N�<�^�������n�̏ ������ڏ�J�8� n�����X�����Ɵ�����SRACFG� �Yk���C�~*�_PARAMSa�3�Yk @���@`3V��2C�`A5�Fby�C3V��BA��*SYS�\�*F`V9.30�146 Т5/2�7/2021 �A��������J�2RED_T �  4$EX_D_RTQ�
��ITP�
�PR�G�
�LINE�*�  �RDCR��A� � $��PX_TORQU�6�  	O�IN�T�THREST� �]�GEAR_R�ATIP\�WARN�_FLGF`$C�OMP_SW-��$v�ER0�SP�C���%�_���J_2TH2Nбհ��� 1  }���PROT_.��_  D �$ENABL�� ���LVL2_PsCTݲ�SEV��~c�L10_CAı���C� � h $�_R�EM~�ST_DATZ�e�^�\�����6!� _�LAi��l\���RO)�%������<��INT��� P �DES�IG6�~��1�1�+Ʋ���10^�_D�SEC~�s��@�F�POS11� wl ��MEN!����б$AT�PERCH	�DO�UT_TYP�Y�INDX��P�'��~�P�TOL~�HO�ME{�P#�2+��1�C�U�g�yߋ� 4#�3+������߸����� H#�4+�+�=�O�a�s��S �&�5+�	��`��������� "�6+�
%�7�I�[�m��� �#�7+����������������8+�1CUgyޝ�SMSK� � $Q�$�EN<���MOTE��� T �1��1�IO� PI� �LOCAL_OP]>uSTART)���POWER� �FLA)��� , }�$DSB_���P��dPC۰���S2327 ��M��� DEVI�CEUSOSPE���^�ITY�O�PBITS�FLOWCONTR� ��TIME� �C�U2 }� �AUXT�ASK���ERF{AC$TATU9 ���SCH�� t� OLD_� C��$FRE�EFROMSIZl���GEj�IR� �	$UPDT_M�=®�PTP	�E�XP�*�#!��FA�ULj�-��RV�k�A�!  �$l�O!  r�VAELk� ]�6N��|1�� �S@�~�	� �$��_$2 ɲGR�OU�r3T��AX�9!r3DSP�6JOGLI`#F4��!b��N �l32�AXʰzi&K� _MIR�1��4P^�TN�8AP� �RPXR	�ʱ����1�ʱPGFBgRKH�!�&NC�0I�  BB�MB�t2P� D6�r3�0B�SOC}63NyEDUMMY164o2SV_CODEz��FSPD_OViRаr���LD�BF�3OR�G� PE�F�)PC�G�0OV�5S�F�JRUN�C��S1FV��3UF`�+Y�TOH$LCHDL}Y�7RECOV�D��0Wi�M�@jU�0��+S�@�_P[�� @��TINVE\�
�OFS�PC/0��FWD�AfT�A�AX��5�@TR���&�E_FDO�6MOB_CM��PBЇBL_/�ba2SV�!��� m�j3�BGg HAMC `� Ne�Rho_M$`b"��L�PT$<�\`�!�T$HBK�!F�a�IO��em�aPPA�j�a�i�d�ese�m�RDVC_DBG�%pA�%pvR� <uޠFx�c<u3Dv�P ��$���j �AU��0LCAB4��ų�P�wS� GhҲO[`UX~FSUBCPU���0Sd�v��S6d� 1��|%c6d��$HW_C� P ��`*��%a� � r��$U�NITVDP�I�A�TTRI� ]��0C3YC®qCA�r�3�FLTR_2_FAI���s��P�;�CHK_� SCT6�3F_I�F_S�܂�e�FS�.bN�CH�Ad�ć�-bW"�RSD�P�fA�#�m�_TKh�up�SM E)M� 2�MJCT
���r�
�%`��DIA�GERAILAC42s�rM@�LOi@б��F5o2PS�2� X,��u�cPR&pSİJ����Cq��	�S�FUN�q!RI�Nx�ı� ���L!RA,�ʰ~��`D�Q��dD����dCBLCURY�u�An�j�q�j�DAT@E���u�n�LD� �@�aף�1N�ܑףTI���m1�r�$CE_RIYA���AF�pP��"��(�T2ĐC��#araOIT��VD�F_L',R�!O L�M0cF��HRDYYO�1�PRGܠH>���1� ��v�MULS�Ef��#�w3M�$�J�JJ�B�G�KFA�N_ALM����W{RN��HARD� $�&� P�"O�2��2!d>�.E_aPFAU� �R�c"TO_SBRmb0j�I�s#����MPINF�Pp_���͡��REG��NV� �>FDxN��TFL;��$M@x�̀�#���`���6�CMpNFt��scON�PI��4��P��P��$�3$YWҶ!4Y2C1���$ �CEaG�r3�@��AR�0M�E27o2�՛� EwAXE�7ROB�:7RED�6WRsPGA_��kCSYD@�ѫ`:�S�WRIsP��)�ST��3d H@�@%EK�� ��8o2B�"�0BM��QT�9˓y`�OTO��� 5�ARY�3��őyt�C �FI)@j#$LI�NKe�GTH���� T_J�Q�D390o2��XYZ�"�����OFF�P���������B�0�`0�vQI � 1�FIx��J�r ��D��4_J!*2�B���a7�c�m�3%a$ [���d����C�EDU�Rr�E3°ړTUR��!X�������X�`��FL��HP�s�� ���P�3�C�Q 1� K�0MD��זp�u��w�#ORQm�H�1J���6ؕ&@O�Ѐ(p��#�1���OVE�W�M� �V� �\��b���!��q�K��AN!���� (�X���05ar�����\��1E)R�1N�	ܒEsP0$蓽Ak��M�<�`h��綡�v��AXvS *2��d�2���%��#) ±#)�@"*א"*� "*@��"*]�"*{�"*1�� "&v�)v�/)v�?)v� O)v�_)v�o)v�)v� �)v��)�!�)��e�%oDEBU!�$�`(Ü�p1�R��AB��ȴa�A�V�` � 
�2MsXѳ5%a�7�� �7�A�7ב�7��7�� �7]�7{�.���(���.1�LABG����*sGRO����!��`B_v��9��CA��g�hF�A��EU��FAND^ �p��q��U��G �a)�J��H��X����NT�jS'PVEL|�Q1Q��9X��Z1�NA?a;���C�2��C��Ӱ]���?�SERVE'Pq�� $$�H�jQ!�PPO��!��P��b�QH�R[p�@л$�RTRQ��
��S���P�W(�2��U���_  ql��qÆERRm���I�`5PQBaTO	QQNL��!$)�Uf�h�G�U%��r���SRE��  �,�Q�U`URA~�a 2 d�b��c �d�P �Q�$� {�X�" ��SOC���P � 4kCOUN�TM� �QFZN�_CFG�Q 4&��ƛ�T�s�bqd3�`Qba �R$qm�  ��0M�ϲX�`'�M���uFA�\#��sX�б{�ykaHW��ѰTq���P�?�SHEL��)r�! 5y�B�_BAS��RSR�����SK����1~g�2@�3@�4�@�5@�6@�7@�8~g�RO\P�a����3NL\���AB�S��n�ACK�6IN�`T_��U7����Љ�_PU��"�	�OU�SP,����sfY�;���TPFWD_KcARGa��6`RE�T⌰P�ཡA�QUE����� ��*"�5�I ���3�s��.�6P����SEM	�Ö�1��An�qSTY߄SO���DI�)�]C����V�_TM��MANsRQ���END��$KEYSWI�TCH.�C�����H}E��BEATMv�PE��LEFbN��@Jt�UB�F��C�S��DO_HOM&�Ol+ӀEF�PR6�POr��:���C��O��<3`�aOV_M��!�E5�OCM�����1��P�P�sHKp�" �D����]pU.b��M���]���FORC���WAR���b�sO}M�� # @z4Tf�T�U@�P��1��В�3��4�A�b�`�OS�Lv�$�b��U�NLO	�,d޴E�D:�  �p�@HD�DN�Q% �PB�LOB   ��SNP9�S*r& �0��ADD]p_q�$SIZ��$V�A�@�eMULTI�P��Õ�Av�?' � $��H¢K��S]C��CB`���FRIF��`S�s���Ƥ�NF�ODBU�P������X�V%�6�IAd�pC�Jtg�XJ�a�q�(� � 9�_bTE�+�R]�SGLK�T�� &?pd�iC�L��STMT)}�PS�EG-�BW� M�S�HOW���BAN��TP��W{�W���h�S	��`V�_Gor;) ]�$PCq@�`��!FBr�P	�S�P��A���`VD���nr*� �'aA00zULᙰS�@��S筰S緰S�5Q�U6Q�7Q�8Q�9Q�AQ�BQ鄰S�;AT愚�S�FQ� �]�1Pj�#����1��1��U1��1��1��1��U1��1��1��1�U1�2P�2]�2j�U2w�2��2��2��U2��2��2��2��U2��2��2��2�U2�3P�3]�3j�U3w�3��3��3�騇P���3��3��3���3��3��3�3��4P�4]�4j�4�w�4��4��4��4���4��4��4��4���4\4��4�4��5P�5]�5j�5�w�5��5��5��5���5��5��5��5���5\5��5�5��6P�6]�6j�6�w�6��6��6��6���6��6��6��6���6\6��6�6��7P�7]�7j�7�w�7d97q97~97��97�97�97��7���7\7��7�7��Y�VPr�U�RQ+��@5�
�pV����Q, x $TCOR|���vaM�P�R	`�pTQ_�`R��PWe�QN�NTS ]C4��5UOV_U��ZQ��YSL|`�P- � 9���:w��.�ਠ����T�VALAU:u��H�"Q�XFwQ�ID_L��UHI��ZId�$FILE1_�d�t$ã�p�uSSA�a. h��@>`E_BLCK�v�Kbf�ThD_CPUdi:�di.�Eso'd�6�YK��R /? � PW�`��l���aLA��S�`��d�a�dRUN�G �e�d�a�dF��eq�d�q�eH��d4p�d�v5�T2H�_LIv��0  ��G_�O��P�P_ED�I��  Lp�pTs1\rԹȀ_a����zp�BC2=�2 ��B�����֡TqFT8˔�tٓTDC�kp��pM���v�q�wTHD��w�	�S�R��<̰5�ERVE̓7��ٓ7�$��q؀� 3X -$b�LEN̓o�ٓb���cRAr��vPW_0Qґc1b��T2��MO$\a�S���I��:R`aщ�Db��DE�����LACE��+SCqC�:R��_MA�p��/��/�TCV6�W��T(�X�w�m�)��"ᛕ�"�J�A�M��|�J�;��)��n�2͠���3����̰JK�V�K�����$��J���7�#�JJ+�JJ3�AAL#�Y�+�Y��S�0�W�5���N1�~���I�3�8TLπ_xy���IrBCCF#��4 `�@GROUP�Pg����N�pCw�~ �REQUIR"����EBU��^���$T�� �_���q�"��t5 \~��xA�PPR�CL8R
u$epNX�CLO�p"h�S�u}��
�qb�6 �`M�p4����겸�_MG
�°C�=�?`̸��1�ͷBR=K˹NOLD˶��RTMOSq�����	JSp�P[��+��@3��w�����6Hŉ7H�Y�3a^��t7�� �����x��+���PATH�ǀ���������è� �6MQ��SCA�r�Y�6��INa�UCՀ��Z!�C+�UM*�Y���`ʐ1��Q=�L�+��L�b�L�PAYLO�A	�J2L�@R_AN�q��L�`�ٓ���٣�̵R_F2LgSHR1���LO���o���.���.�ACRL_�����ԁ�9H�P8R$H̲?�FLEX[�ġJ�v8 PE���6��H�2b\�a�9 :n�������䃏��0�������F1��6� J���я�����z�E#�5�G�Y�k�}��� ����Qn��̓�^�@�ԟ�������T�OXWQȑ������ ��"�4�F�X�\�e��S�w���������04[�ɤ: ��p֯�����@ATc����CEL��Eq5#�J ��9�JE��CTR��^�TN�A1&�H�AND_VB8R�[��P��; $� Fi2̶��SSW[������<� $$M�й�P��(���, �%6�6A�P�м���Q-9ŽAּ�P�A���A�80׻}`�D*��D�P��G�`�9CST��1���1N�DY�`V�̶4@5�� c��������ц����� �PP�Y�b�k��t�}ņŏ���u=1 � ��� ���E<���AASYM��ZP	���<<Q����_3p�&�9�#�%T�( C�U�g�yߋ�J��C����S�Y��p�_VI�#h��`V_UANsr `'cH��J� ?bmE?b��Cd��Pdtf ��C�$�6��e aL�T�"�pHR�p��q>�"�an�hrD	I� �Ot���`ɣ�? XG2I*QA G���Aqd�OSOsg�A ��e��` @ �� �!ME��Мjr�bQQTpPT@�P����q����G���P�x�q�yT�P��� $DUMMY}1b�$PS_a�RF#�  ���vn��FLAˠYP����s$GLB_T� 
u"��pv���b!nqA XE�����STđ�SBR���M21_V�T�$SV_ER��O�|Ph���CL<�h�A���ODr�`GL	`E�W̡B 4Ӡ�q+$Y�Z�W˃���Ѷ#Akp*�VRD���U��C � N�倭P$GIr {}$�� B��8���̡D LӠ��{R}$F{RE�NWEAR��Nh�FU����TANCh�eqJ�OG�9� E � $JOIN�T��  ��MS�ET̡F  �E;�e��S"���̡_G�  j U���?��LOCK_�FO���!pBGL�Ve#GL��TES�T_XM[���EM�P���#�:��c$U�ం2C���I�D�� �I�B�j�CE���j� $�KARMsTP�DRA����~�VE�C������IUI�E�N�HE�TOOL�*�V)�RE��I�S3��ݢ6k�^�ASCH�� �FʡO�Ԛs�t3���SI�K�  @$RAIL_BOXE���ROBO�?����HOWWAR�G�9��p�ROLM �r_���p��'�R�n��O_F�!���HTML5	q�%%� #AC�������H���R��O��I`��"𓑗��OU��'J t��E�BQQ;"X!��PO�B PIP�N� Ӣ'����p�I�ʰ��COR�DED����R�X�T8�	�)��`�O�Qp K D !�OBm1?#Ǉ���s ���{PA!SYS���ADR@!�`�pT�CH�  L ,�� EN�bw�A��_�����[��VW�VAmqM � �����
uPREV�_RTzA$ED�IT9�VSHWRB�T�Xб�Ł`�D|p@o�H$HEAD�Q�`�МQ�A�KEŁ�pCPwSPD��JMP��=L	uS�TR��,t�N��l���I$�S@"C� NEƠA!|'OTICK*�QMu��fq��HNJ�O� @�������_GqP7��x�STY���LO<�����3���P�
4�G��%�$��=T�S6!$5a�q�>p�9PP7�SQU���<� aTERC�p�z� S�Q ��`��� ����B O�p�sl�IZ����qPRj��qU�����PU!e�_DO�Z���XS��K	vA�XI����N�UR  ��A"@�%�Ʊ! Y_����ET��P������E��F�G��A�AQ�t9�2�X��A�SR�$Rl��)��*@�& R	2@7@)9@99 �[7�k7�{6�� �9���B�	C��C�t_�_�_�T��S�SC$��� h��D1SE����pSP;p�ATi02f�$���~�rADDRESǣ=BD�SHIF��@��_2CH@ ��I\C�!�TUC�I�!� T�CUST�O����VԒI/rU�����I��@
#�
�"V�u�opV \R�����T,#����"C�3&���c*Ɔ��!��TXSCREE��Wp��TIN!A����$�����@X T�у�I� ����_�16����-4@�RROD@o������*1���UE���Y ��@���pS�����RSM$���U`s���	v�1�`S_ރ��6.S�1�9�7.S��Cx䒗24 2X&pUE�DZ5r���6U�WGMT�`Laa���o�/����BBL�_�W�pop[ ��` [BO؁gBLE��rC?�*"qDRIG�H{CBRD���C'KGR�p�ETt��G>�AWIDTH�e�����ǡ�U�I��EY��nq\ Ad����^�g�'�Q�BACKe��rU���upFOa�)WLA-Bp?(upI�蒏$URE�VPAI�_{pHQ1 ] 	8�ao�_��"yR|pRŀ���q  fQ)O�op^.����@�U�@�SR��j�LUqM�S���ERV"�����@PY��D_sp��GEZR@���zГLPe��E����)�6g��Dh�Dh�Ci5*Ak6Ak7Ak8&b��@2�P�Y��$�v���S��^�AUSR���` <R�{pU�
�9#
�FO' 
�P�RIm�3�pT�RIP#�m�U�NDO��a� ��1p��Q����@A������ btR�`T�G ��T��e!orOS�q�vR��W2[sáAc��̃ӎ�rG�$�QA�U!aAd��p�3!bF�[sOFF�*��e��sO:�J��c�$�L�d�GU��PK���g�bq�Q�SUBG� ��E/_EXE��V��[s�WO[ f�p�{w��WAD��`��z>P�V_DBŃ�݀+rSRT�p'g0.�n���4�OR��'RAU9 �T#���r�_7���h |B ���OWN^p��$GSRCb0�0��D�<y�7MPFI^���ESPa�,�� ե��S��W�E�R�Ai# `�p����"���7COP�$G�`p�_������ςC�T�C�������  D�CS]�P�j4ζCOM�`{@ ����'G���sہ�#�6��VT�q*�pv�Y��Z�
�`���l@S1O#SB��P֨
�40��_��M�Ü�5�DIC����A�Yo3�PEE�@T�[Q+�VR	Л��!$�� 9�vP۠(�ԡ >�R��>� �wͤ�p���L�:# k$2?SHADOW���~��_UNSCAI�毳OW���DGD}E�LEGAC��I'��G�"l ("@NO�P�TY�&�L���VW���G��Am � ��VqEb3��<�ANG�4�J��J��s<�8�_X �w��w�b�|�q��3`�$p O���VF����VCC����n7�C��RA�����΢: A�$��_^�� l#pG�{@mN��`|��� STEգ���P� ���P���pH@�����p8O�}���P_A�������h ��Ao� N�O� ��Y��þ����S<`C
`��DR�I>���/�V@���B�U��s��MY_UBY�d�ͫs����� � ��N�ȣ�A_��k��n�Lk�BMnA$n�DEY|�EXyќ���MUL��U�Mư0USHq��p_R��!5�p A�G� PACI��,���C��@���s��3h�E�R���qt������pS $ ��G0�P�"HF�Ӑ��R�p��q�@��PP1�A��	�AX�0T�SW����v��2��SGA�BA����@E�`UEe� YQ@��HK�rr�P���G�8 ��60E�EAN	��
���0���MRCVAs ��`O��M
��>P	pJ$�C�JREFGG�lS>m�A��N �`O
�`
�q�S��_v�
�'��R��n4��r�4Dt ��� ����a�y�COU}�p���,�o\�ƀ2p"@� � 	�pqS"���0�+UL7�rƐC=��Q3s��NT����ϒ��Q��a��L ��%ȣ%�Q#'�a��wTCC��u t�p3MD����HU�H�vc$SAD�CMP�aFi&�%z%j _Dp�AR�ĝ��!"X�)�l�GFL�3v,+ &Z�%#�_`0���%�o�RO�@92��D��P��P��URE�RN6��RI��l#INрuJ�\�nˁ���X����IN��Ha4���@Vu���L��3�C�5WU�4��������:I��LOo���ܱD8D�iA�aNSIy����� ��F��F��X_�PE�8Y�KZ_M$Ӈ�W3@���Ä r�KR�G�#RSL<�'w �t1��M'p�b)g=y�C��G�Q=� ����s�"�f >��/??(?���c|`l�f�` PIA��wx ���HDRȀ���JO�`t��$Z_UP}�	�_LOW>ea�� ��LIN�rEP��s|y.aa���p�Ɩ�a�����y� 5�PATHz*p �CACHpD ]A�e\AP@�i�����C��IسF6�tT8E�t4$HO
�l��`[��Ӭ��S=v]x]���PAGEaƞ�VP@򭠊r_SIZӔtZ���x}Ә�uρ��MP�z�IkMG�[@AD�y��MRE`��wG�P]К����ASY�NBUF��RTD�6�B��qG�LE_2�D��^�BBPC4�U��\@Q��&�ECCU3�VEM�e��wVIRC�qV�>�ૢB�3@��&NFO{UN�DIAGR�Ry�XYZ�0����Ww���1����`RT���IM��U�ނ|��eGRABB(\Ԥ��LER��C�b�F�"�a�V50�������ϑ �eKz� Z�BACKL�AS�`��aX��{�  �s�TA � @�?�7�$�a(���| A��1� ǂ�3'�T�� � �ї`�R0�IN�4�t�`B��EVEц�PK����]G�I�NO�a䱽�_�HO� ��} � �]���l#�0`�˦S�H`��ROD�AC�CEL�P����VR�U�`l����Ұ6x�AR�PA�.���D�REM_Bvה �_JM�@�x�~��%$SS�C9��q�\@���� �@\AS�WFNܵ���LEX�� =Tj ENABi@&���`�FLDRA�F�I`�B��A؊� �'��VP2�f�'� v1.pVl$� MV_PI��PĚt �0U���w0j�Fh`��Zqʍą�T��1vȚ1̅�C�GA��� LO9O�S�JCB��Y�΄sCON�po�PLCAN=�tҢ�!F}�Ưة�p7�M^� ��]�f�S�P�+�}њ1�+չ��1R���Қt����RK�B)�VAsNC㳽�R_O� T�� (j �C�C�3 �3vRV0��A��T�� 4_ �����0k�8�e�x� h��}�8a�mFOFF~��a�;�S ��dEAwY
���SK
tM�V�VIE�2� ���p�R� < !ݺ/tdI!��W�' D��e�CU�ST�"U� � �$�TITQ�$PR��C5OPT<Ð�q�VSFQ ���R`mF[8O�K�MOT%���޳&��J�*M ZDO��� D��_aAL�I�M}p^bo�I��$_MSG_QV�O�H�t� �q_�b �����3�� g`�Sڀ�X�SU$� x)`MSGPD_��_aB�P@	�SA@NB^bLNTKcMPKd;�C�`��&�a��4Ų��XVRU#��ϒ3�T� �Z�ABCJ� xѐ�/s  
! �����VSp` � � ���df�IV�ځIOmB�$Kv�aITV�sT�RGTDV��
0J�����pDI$`�� K0�P�V2pځ�PZ�ځLST��ځA R�A�_ST��|e���DCSCHW"G� L��dOa��scg@A:pSIGN�� ���ځ�_FUqN8@ڀH�ZIPT$S���u�LDL��� y�ZMPCF���Y�E c�qX!D�MY_LN�����D!EP�� �$IqL0]$CMCM�8PC�sC�A�!4P~� $J�#�$Dq�"�"�'rp�%�rp�'_G��R�"�'U�X!�\%UXEUL 8!��%5�%1(1:9x(1J7� FTFL�&�w4ޑ�Z%�������� Yg`D�p� � 8 �$R�pU�$H�EIGH�3�?(�z� ��Pƕ�� �àA�L1� $B�X``��k�_SH�IFcC��RV��FL@p� 	$5B�C%` �"�Ap�A�W� ��'�dxCA�D�H�CE@ )V� P9PH�Q�� ,z��8�?�9��$RBTIF �ϐ�������A�@CVT�b��C�AT��@D�CR�R1�A�A�5`� 	� 8��2�AE�ĳ��AA�T��S^XGP�A���A����A��w7b_�_^_ ;����;`H�;�S��;�d�;��Y;��*�_pv`�_ o�] o 7oIo[omoo�o�o�o��o�o�o�oS(QIO&�� 5US�_gRED�Z5W�@P�TBH�SE�Sy/Q2e{ �FQB�xp��z�_���_��(���Y�%�6���hW5U������ я�������)�O� o�t��E;��������� �ӟ����	�?�a�f� ����!��������ϯ ��)�K�P�o�!��� �����˿��ۿ�� %�G�L�k�-��mϣ� ���ϵ������1�6� H��i�ߍ�{ߝߟ� �������-�2�Q�� e�S��w����������=�.��CUwINGT 2���Q�q�FQG;� l�~��r�_<��gXf�0 ���� ������P> tZ������ ��(L:p� h����� /� $//H/6/l/~/d/�/ �/�/�/�/�/�/ ??�D?V;UqFPOS1� 1$y  x���qs���?�? �?�8�?�?�?2OOVO �?zOO�O9O�O�OoO �O�O_�O@_R_�O�O 9_�_�_�_Y_�_}_o �_o<o�_`o�_�oo �o�oUogo�o�o& �oJ�on	k�? �c���"��� 	�j�U���)���M�֏ q�ӏ���0�ˏT�� x���%�7�q�ҟ���� �����>�ٟ;�t�� ��3���W��򯍯�� ٯ:�%�^�������� A���ܿw� ϛ�$Ͽ� H�Z����AϢύ��� a��υ�ߩ��D��� h�ߌ�'߰���]�o� ��
���.���R���v� �s��G���k���� �*������r�]��� 1���U���y����� 8��\����-? y����"�F��C|h52 1t?0j��/ 0/�T/�Q/�/%/ �/I/�/m/�/�/�/�/ �/P?;?t??�?3?�? W?�?�?�?O�?:O�? ^O�?OOWO�O�O�O wO _�O$_�O!_Z_�O ~__�_=_�_a_s_�_ �_ ooDo�_hoo�o 'o�o�o]o�o�o
�o .�o�o�o'�s� G�k���*�� N��r����1�C�U� ����ۏ���8�ӏ\� ��Y���-���Q�ڟu� ����������X�C�|� ���;�į_������� ���B�ݯf���%� _�������ϣ�,� ǿ)�b�����!Ϫ�E� ��i�{ύ���(��L� ��p�ߔ�/ߑ���e� �߉���6������� /��{��O���s��� ����2���V���z��x����3 1� K�]��� 9?�] ���~�R�v ��#���} h�<�`��� /�C/�g//�/&/ 8/J/�/�/�/	?�/-? �/Q?�/N?�?"?�?F? �?j?�?�?�?�?�?MO 8OqOO�O0O�OTO�O �O�O_�O7_�O[_�O __T_�_�_�_t_�_ �_!o�_oWo�_{oo �o:o�o^opo�o�o A�oe �$� �Z�~��+�� ��$���p���D�͏ h�񏌏�'�K�� o�
���.�@�R���� ؟���5�ПY���V� ��*���N�ׯr����� ������U�@�y���� 8���\�������϶� ?�ڿc����"�\Ͻ� ����|�ߠ�)���&� _��σ�ߧ�B��߱���4 1��xߊ� ��B�-�f�lߊ�%�� I��������,��� P������I������� i�������L�� p�/�Sew ��6�Z�~ {�O�s��  /���/z/e/�/ 9/�/]/�/�/�/?�/ @?�/d?�/�?#?5?G? �?�?�?O�?*O�?NO �?KO�OO�OCO�OgO �O�O�O�O�OJ_5_n_ 	_�_-_�_Q_�_�_�_ o�_4o�_Xo�_oo Qo�o�o�oqo�o�o �oT�ox�7 �[m���>� �b����!�����W� ��{����(�ÏՏ� !���m���A�ʟe�� ���$���H��l�� ��+�=�O����կ� ��2�ͯV��S���'����K�Կo�������5 1	�ߥ����o� Zϓϙ���R���v��� ߬�5���Y���}�� *�<�v������ߖ�� ��C���@�y���8� ��\��������?� *�c����"���F��� ��|���)��M�� ��F���f� ��I�m �,�Pbt�/ �3/�W/�{//x/ �/L/�/p/�/�/?�/ �/�/?w?b?�?6?�? Z?�?~?�?O�?=O�? aO�?�O O2ODO~O�O �O_�O'_�OK_�OH_ �__�_@_�_d_�_�_ �_�_�_Go2okoo�o *o�oNo�o�o�o�o 1�oU�oN� ��n����� Q��u����4���X� j�|�����;�֏_� ���������T�ݟx�����%���6 1
(�ҟ�������� Ɵ������>�ٯ b�����!���E�W�i� ����(�ÿL��p� �mϦ�A���e��ω� ߭Ͽ����l�Wߐ� +ߴ�O���s����� 2���V���z��'�9� s����������@� ��=�v����5���Y� ��}�������<'` ����C��y �&�J��	 C���c��/ �/F/�j//�/)/ �/M/_/q/�/?�/0? �/T?�/x??u?�?I? �?m?�?�?O�?�?�? OtO_O�O3O�OWO�O {O�O_�O:_�O^_�O �__/_A_{_�_�_ o �_$o�_Ho�_Eo~oo �o=o�oao�o�o�o�o �oD/h�'� K���
��.��xR�8�J�7 1U� ��K�ɏ����� ��5�Џ2�k����*� ��N�ןr�����П1� �U��y����8��� ӯn��������?�گ ���8�������X�� |�Ϡ��;�ֿ_��� ��ϧ�B�T�fϠ�� ��%���I���m��j� ��>���b��߆��� �����i�T��(�� L���p������/��� S���w��$�6�p��� ��������=��: s�2�V�z ���9$]�� �@��v�� #/�G/��/@/�/ �/�/`/�/�/?�/
? C?�/g??�?&?�?J? \?n?�?	O�?-O�?QO �?uOOrO�OFO�OjO �O�O_�O�O�O_q_ \_�_0_�_T_�_x_�_ o�_7o�_[o�_oe�w�8 1��,o>o xo�o�o o>�ob �o_�3�W�{ �����^�I��� ���A�ʏe�Ǐ ��� $���H��l���+� e�Ɵ��Ʂ����2� ͟/�h����'���K� ԯo�����ͯ.��R� �v����5���пk� ����ϳ�<�׿��� 5ϖρϺ�U���y�� ����8���\��π�� ��?�Q�cߝ�����"� ��F���j��g��;� ��_���������� �f�Q���%���I��� m�����,��P�� t!3m��� ��:�7p �/�S�w�� �6/!/Z/�~//�/ =/�/�/s/�/�/ ?�/ D?�/�/?=?�?�?�? ]?�?�?
O�?O@O�?�dO�?�O#O�O�o�dM�ASK 1�k�B�O�G�GXNO�  �O�O^MO�TE  \  �QU_CFG �\^�T�jPL_RA�NGXQTA�e��VO�WER �e��P�VSM_DRY�PRG %�i��%YO	o�UTART� V�VjUME_PRO�_�_so�d�_EXEC_EN�B  �D�YG�SPDL`�`�hΣhTDB�o�jRM��o�hIA_OPTgION�TiQ�S�lQINGVERS�q Zbo�II_AIRPUR�P� Tj-T��KMT�_�@T�PZ[�UOB�OT_ISOLC�\��p�q�]�rNA�ME:|�J�|_C�ATEGX�S.S�%PU�]�0�ORD_�NUM ?�X��qH727  �D�������@�PC_TIMEO�UT�_ x�@S2�32uR1 U�c� LTEAC�H PENDAN�܀qG�U�P�L�XOV@Maint�enance C�onsRB(��F"�D�RDNo Use8�t�:�������Ο8���B�NPO&`ނ�Q$u�CH_eLO`u|�D	c�~.�!UD1:��z0�R�@VAILy��u�UlQSR + v{"q�Z<��R_INTVAL�v��Y�~۩V�_DATA_GR�P 2 UiQ� D��P�O���O ���� Uοܷƿ���  ��D�2�T�V�hϞ� ���ϰ�����
���� @�.�d�R߈�v߬ߚ� �߾������*��N� <�r�`������� ������$�&�8�n� \��������������� ��4"XF|j ������� B0Rxf�$Q��$SAF_DO_PULSYP]�U@<�Sk�SCANՂv��V��P"��"6��a�U@U@
��U@!��s�s�!RB ��N/`/r/�/�/ �/7/�/�/�/??&?V!�-��"2O4�!Z9dO8LQnU@��
 @�[�?�?�?�8���P�5��_ �0RBT"pwCO�/OAOSOED�� ZO�O�O�O�O�O�O�O __%_7_I_[_m__`�_�_����9~=��_�_�A$�;�#o��"a�qp�$��
�u��Di��!&!��� � ��vA&!�!��! "a�o�o�o�o�o�o %7I[m� �������!� 3�E�W�i�{������� ÏՏ�����/�A�S�e���?�������� ҟ�����i�<6G� Y�k�}�������ůׯ��*��R0�2tcBe ~o;�M�_�q������� ��˿ݿ���%�7� I�[�m�ϑϣϵ��� �������!�3�E�W� i�{ߍߟ߱������� ���v�/�A�S�e�w� �������<���� �+�=�O�a�s����6ta��`���L0����� � �!�������� �c,>Pbt�� �����( :L^p���� ��� //$/6/H/ Z/l/~/�/ej�_jB�/ �/�/�/? ?2?D?V? h?z?�?�?�?�?�?�?��?	j�/O<O	f����b5Om	�12345678�[bh!B!���%`*��Q�  !�O�O�O�O�O__ *_<_BQ�/e_w_�_�_ �_�_�_�_�_oo+o =oOoaoso�oqMT_�o �o�o�o%7I [m������oBH��$�6� H�Z�l�~�������Ə�؏���� �2��k;!7�>�h�z����� ��ԟ���
��.��@�R�d�v����iD� ����̯ޯ���&� 8�J�\�n��������� ȿڿ�o���"�4�F� X�j�|ώϠϲ����� ������0��T�f� xߊߜ߮��������� ��,�>�P�b�t�� Eߪ���������� (�:�L�^�p�������������qD�F�����6HZvJC� �A��*   ���(2�" _}�h
�-V�	�.B2�����h�/%���@1� 3 4 5 6 	$z�� �����
//./ @/R/d/v/�/�/�/�/*M��"(�"P�/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO0OBOh0%���<wD mE�  ��K�OUF��B��t  Ў �I�OUH`2�$�SCR_GRP �1"Y�"�b� � �2� �	 � "P5QER>T&fCU_@UGQW_m_�_3@��EP�� �RD�` D�@:KS�P� �Q��[HR-20�00iC/210�L 567890r� e� RC%`�)`0
V09.01 T`tX�Q6�A� xf4QUF#Q �S#QHvA�QBW��k	zb�o�o�o~UL��H�g�5Z#R2H�á�D�X��Bo���f\������۟�BE��a�� 6�n �J���3B�[�@BXzR��WߩĴ�'UM:��>udp�hpjlp�g�2�_��_�T]H�{(ohj@�pY�B���B�ff?B�  B�^�Y�Gƙ�\�m�PQA� �|��P�Q��PQ�Q��  ?���P�| ̏���PQF@ F�` �����#��G�2�W� }�h�����şH���Ă`�۟����B�� ��e�P���t������� �ί��+��O�a�@G�S�_����`I
���׿�T�P@��A�Ed�\ń����B�~2�1234(c>Ǖ��mϮ�,Q@�ýuSP��H�2 �����Ϯ��� ��.����+`�r߄� G��ߓ��߮�
oN���	�c�PECL�VL  2����b��+v�L_DEFAULT$���3~8�HOTSTRD����X�MIPOWEKRF#�rP�z�oWFDOE� P��QERVENT �1+�+�q� L�!DUM_EI��/���j!AF�_INED�	���!'FT�﮾��\�1!Wvx����K����!RPC_MAIN�����������'VIS�������@!OPCUAA殺/�!TMP PU���d{��!
PMON_�PROXY���e �$����fp�!RDM_SR�Vq��g_�!�RP����h�/!%
��M;��i�T/!RLSYN9`�p/��8C/�/!gROS�﮼�4�/��/!
CE� MT'COM�/��k�/8?{!	2CONS9?���l'?�?!2WOASRC���ms?v�?!2USB�?���n�?O!STM��6O��oOhOo���OYO����ICE�_KL ?%��� (%SVCPGRG1�O���E2�OD_�@3%_*_�@4M_DR_�@5u_z_�@6�_�_�@7�_�_�@���_�A9ok�D�Bo �A�Ojo�A_�o�A?_ �o�Ag_�o�A�_
�A �_2�A�_Z�Ao� �A/o�QXo�Q�o �Q�o"�Q�oJ�Q �or�Q ��QH Qp�Q��Q� :�<Q��O�B�@�O�@ ��ʟ�Ο�ݟ�� :�%�^�I�������� ��ܯǯ ��$��6� Z�E�~�i�����ƿ�� ���� ��D�/�h� Sό�wϞ��ϭ����� 
���.��R�d�O߈� s߬ߗ��߻�������*��N��J_DEV� ���M�C:Y�k�GRP �2����@bx� 	� 
 ,*����Ւ����b����V�� V� ����,��P�7�t� ��m��������������(L^���J�໒�c���� ������0 B)fM�q��@���//qo��r�����C/Q//�/ �/�/�/�/�/�/?? B?T?;?x?_?�?�?�?D�?)/����?O 5O��YO@O}OdO�?�O �?�O�O�O_�O1__@U_g_N_�_�?�ಒ�% ���_jN�_�� s_�OooBo)ofoMo _o�o�o�o�o�o�o�o >Ps	��� O�lO:o�r�� #�
�3�Y�@�}�d��������׏���������=�tD?�{O폆� m��������ǟ�� ��:�!�^�p�W���{� ��ʯ��������� ?�Q�8�u�\������� Ͽ���ڿ�)��M� 4�qσ�گ��^Ϸ��� �����%�7��[�B� ߑ�xߵߜ�����������3�C�d �Tߚ6�P	 ���������$������ͭ:����QC�a�?�R����{	@�d����Ơ@-#�@Q�����A��A�cN��Ը�B�EB�oz��ۃ���'��v��-A�<��A��A���&�1k��Q�%�NORMALIZ�E_HEIGHT|C�N�T�@�\��`�=�l���|�=E���'���=���к;�	����T�`��ja�����@����?�D3@�t�����>��h�T�A�1B��9�}�����B��jB�E�c�I4�T�?G��r����A`�8�@xh=A�?��@�!dQ�T��%	� POFF�_APROACH��*�Q�6 &�`�D�#����Z�/�K?0D��A	u��vO����`�@��g��A@=�`����
@�%��R�Z(
2�?B�U���Qt�����BBOB��G�In3T������B����;�A��	����������RS>J��G�Ꝙ�Q�8�>J4�@�����9��R��ք�{���A9�����S�X@թ�ﾌ��(
����BU���S?`��ו�BK���B���tr�����B�5��N9�A�{��I����*����\�=�\��<ؑy=����=W����ȳ�<�S���J�����@s��O��*�@ss����
>}�|��A�c�o��E���B�,B�]�2� �T�=��q�����A?��@�A���V@u�p�JOGGING �ATION�j(Tכ�5��V�5=a��<���q���B;�4������#��f@h����@�z{�Ϟ�>�!���A�~���7�D,��B���B�g��/. ���A\���@h �A��@�"�D/V!��l/��9�=�	��=�L==�tD���J<�V���Β� bn@�F��@o"��%�>���(
�_��A�ː����D)zB��s�B�f�� �� ����tAI�'E@l��A�?�@�@2?V/�Oz"�\�А��=��>YQ���P-��qW�=4�w$?�����-�@�[�|@	��@j�?+����>�0(
��
�AהO���#��C�RB��lBˏ9�>�����A�uq�@��yA���@���?�*3LOo-�\�>�
�=�q%>B�H�=� l��?a�<O#������$�Q@������0@��~���PÜ>���Aڰpk|��C�B���B�/��-�- ��
Az��@���A��B?�״��O*3FE_�21�Os)���D��= k�=ե�=l� �*;�y�T��$�@��W����@�X����_�>��q�Aލ������C"�B��B���� � *d~P	&7A�~��@��A���@Y���_�*?�oz"Ŭ�w��=�c�>:��=���c���<D����1'��_@��߿�0@��U[���Q>����H[D�A��c��C��'B�QnB���/~P�A���w@�A��L@z8ho��1Q�o�\��/H>�>��1U��3�����=UǇHN��2��+��@��%C@J$l@}�����{x�@�ւ]A�7����l;�B�B���B�j@m���� �A���@Y�0A�?��@�w(<N�3�z!���϶�=f^=��2�=R�R�]�$����&m�&@��߿�+�@� ���>(
���{BǸ���`�CO8B�,tB�p�}�?��{����A�?0@ʵ��A�`i@U����"��F��xv8��l>�,�>�&���\格�>_x=����?y���-{@�!|�@6Β@R\��ɔB>��(
���WB_��Z��D�1B�?�#B�q}�r��A�y�@���A��M@������?۟z!�xvG&#>�`��>��$�eP�-�=���uP�?�1]Ae�9q��@\�G��h����SBF���}d���B�2?�B���~Qa�LA�*�@����A�Y�@����ʟ���t(F!�ԑ<�CR=k�]��T �l?*<Ts�HN�!�(�@�V�M�_e@U�U�r�N��`�B����}�h�E,B��0B� @m�>}Q%�A���L@�4A�}��@�ۭ����R�O��n-�(F���=�H�>AH� ���r�N���=!����p'�̭@���o� �d�>���BV���z:��E��BB�fB��l~P"��A���@��A�?8�@b}�`�zcؤ�|�r)	(Fr���=��!=���Ľg�D�	ß,<�|���p,�1�@��4@/ܚ����Q�>����B ݪ�tF���G'�B�ԟ�B޿d�~P#���A��^@��e�A�9V@9C��4�zo+�j�(F�{�=�w�>�;l��o���'Hm=q0��0&��t@�e�@&��`���CpN��sYB#�U�q��5�G2 B�?ۅB߮�l_~P�+5A���@�P�A���8��O��f�<(F�g��>(�>����I
��8��=� h@�a%��<@�Z�0�x����H��>�_��B(xo�n��7�G�jB����B�'�����-aA�;�@�יCA���@��m�����z��b�xv_6�>����?&(���y���.��>p|HN��+�C@�`�@$Y�@v����(m���X��B*���l�9��H2�B����B��7����1%���A±�@ޡ����/�I�CK���(F�;��>c�p>�D�d�������=����H⁁߹�@�N��c��^��n���B/|D�iq���I3�B�w�B�r\��0)���A� LA;]��2h�l������
�
#(F�m��>+ȹ>�ݾ��ߴz���,�=S���h0��"�-@�pP�@��@G�q���{����ś�B4\��e�D��J��B��b�B��'��Y0���A�A��A�����K��L��3�l>��w?�?�W�J��Cr=������`�vJ�@���@��`��m&����B6��d���K{B����B��M����r��2s�A����A��2JÄ<,r�LEAV�_�{(F�`���u�w_����@���B����@���@A�@�S�X����B�9w��b$��L�B��~B����0�0/�g�Aȱ*AKvA�7%0�:�/^���V���>I1��>�m�=�����y[<����^�7���@�0�m @���d�� �>}��:���BAO���\U��Nv�RB�L#B�=�弎��0= JA����A��Au�3@�	;�/��/�?����r���>�%�!dA���ҧ=�J�@�R�b@�m@�,N0a�<�����h��>IBD���ZU7�O�B�cIB�P��>�q>��A�t�A
٩ ҇�"��?�?�O����֐>i��{>� þJww��^ХP[��Y�L�zH1�@ P��ف�����X�BF���Y&d�O��B��B�$#���#�:C�A�tA!�,��(	|O�Os_�B�1�Ql>$��>�7O���Ǽv=u���N��`@��l�@��@y�����&n��[wBH�;�V���PŽB�?��B�O(�R`�<��AگdA�9^A�a�@�O�P_��Go�BX���&]H>�%��?%��b����bh> �|�����@���l(�fD3�����h���#BLz��T�x�QG��B���B��π?n�@^=A���^A�A�C���^_�Fv���*G>�+m>�ڦ�!~��\� O"��R������B��`��>���ьޖX�BO|��R��/�REQB�&_�B�ͼ����?xcA�_�A��A��%@�W���o���B����[#>o���>��������r`��"���<�@�wA�@#x�@PK_���a�侕ǡ�BRK��P�>��S<�B�V��B�6��V*���C��A��&�b��j@�����
Ï�B�6����>2�p>�<�+=(? �����,?>0��oY�@�^�3J��@���5��-�wBU���Nu���T]7B����B��J(_:PC��A�r�@���bAxɖ@��⠏6aY_ER�ROR_MOVE�_��GRAM�N���cfG>W��>SN۽Sݎݻ��ʐ�>(��ҧ�Q?�4�P@���5���]�B[���J<b��U�dB}�a�B���P@�k��4�I�?A�?�AJ���)�3oh��
6���>T98>���)=N�`�����=#Rx0>��)���O@�������@�t]���W,N��B�^6&�H����V�hB|�VB��
-�.����L�3A�KKA���Am�@��ǒH�Z�?�~�6�6u�=0v��=�O�<�U��Τ�<�M���v��D�2@�޿r��@v����{侏 �Ba��}�FD[�W���Bz��B�E��^>�U=�M���A�rEAU��Ay�@�����.��~��5>�G&#>���?�:��=��3�V��=��#0>��Z}��~3@�� ����@����4��z��Bie��Aq���Y�pBw'��B�һ�.��R���A���A��qA_�2?�Ð������ h�,���=�|�>NL�>E7���l]<��S�x��� �
�@V6P��T�@��o�����>���ڊ��A��"!&��5��zB��[BÿZ�Ǒ]�`�9��W��RvAT�9�@���A�C]}D���x������`�G>1!�>��?��YyA�#��=�i������ �@t���@h�@n-?$�É�>�Pd����A�D�������5��B��8�B�&�בz94:+ڰJ��A_Lz@�g�@���]���ð����!�6V����X潄�?=��;�*�W�������@�����$<�,A@�Wߵ=��>8����A� �k��6v�B��nB��]�D�?���e#A�ػ@���Ae��0��l�jc���"&��f0�=kH��=��Ľ�Y���qW<�s���neq.�@�>�|D�K�h�I0>�up
b�A���*uk�7B�uB�4
B�l�]D�<̺a=�A�3@��!�A��@����S?AFE_32f�o��F6JI�=��=�������v�<
�m�����(��@��_��������\ӇB�p��e��7�B���B���DD�B��%A��@���HRd����v��6�#<���y=���<��(����;������$:��@�C���u5���=�Z<L�{�Bb��%��:�lB�/˯B؈�D�AJ����!dFA�x��@��A�@�hg���, 1�4��#�6�H�G>'py>����=�o���	��<��x�������@�=޿�9�@lk'����B>R�Z�*6i��B4���h����A:�B�h_B�XR��^��1�0��e�A��@�]���ϳ/
1$76����>(�>�c�)=U������<��w�������@ʭ�{\�@i�����>DJ�,+'B?��ap��D�$B���B��v�D�@J����=�$A����A��At8�y@=��LEAV����(��+��=[�=�=�
<�?���(l����7�V @Ԑz�k�)�R��0�%�BJ�4�Y�~�GJ�.B��7B��ʔ�=s7A��M�@���A�?<B@țOd?&�93�?��&��@��N��$��@��@������͠p�}���l@��٘��&v@�a�<@�Z�>��քY�þ��Ao{����Bn�aB����B�������Y�����hA����$
�A�?ʯ�lu8O�Ϭ/_�Q|#�鄲��u?���@��j���U�+��?>���?����Z���)�r�@�
@.��@�I����_D��`�YA����P"�Ot@��:�BL�<B�q��&m��Z� ���F�8A���0��oA��/�
JZ�UF_RIVE�TLOC�/iT�5�6 &���[l��^J���b��>��:>�d�N?��ja����A�"��@����	����P>�����iB'���s\bB,���B��B�?��I4�̺�����hLA����P�A�cU�@�ۭZ	NO?RMALIZ�TO��gT�;�f���H=^J=��2ӽk�f��?�=<I�9��fp��@���?�ͨe@U�U���O�=I�A�M�}B6a�k���A��yBr��B�		�In]3̾7�*�!�Y1�&@�ןZ�VIS�R�_�|�T�N�e>s������f�7��N=�{0=�<i�]�;z������AC�T���@��I5>����(����B:����c��B���Bp/�B�s�`}@������A��p���r\A�a$@J�ÄZPLCHANDSHAK"_��lQ�vc�����@��;(=wP l�09<T���h���~�A#!}|���/Ơ�� �8~k�B<����bÒA����Bkr4B����4�5B��������A���@O�\�n���js�|��Ƒ>���>�'}��g�D�&Z��?����Z���<@�+�?�J�@��>���=�����B�W6��P��B�V;cBx4�B�j�}`ڰB�W�A���y�N�b��_&1U���vk�L�=��=�^��)~��>x��u�Kb�	
u@��3?���1@���Q=(����?�BO,��V���B5�4Bn���B}K�4�5Щ���r�C�������Q��U�3	�;�&2 M�3���,�]xl>�hd�?].>�L�����G��������bo 2�H���*��@j�?+@�pP=i����)�BK�e��X�,B5��Bp�5B~�&���?��{P2������1�A��L��ǒد�/Ͽ:���,�e$������:�=���>��=����N0���P�A0��t�]`�������Em<�����oBM��W�]�B51 Bo�BB}�O��G��r��^B�����<FA�3�ߔ��LLҿ��ם@q������{S|>��w�@��T�Z�,�>�;1AQɛ��J�������@�3���`��@۸I��l���m������L�x@�¼�'B��B�ߓIǡ�;{%�����A����AP�{A�OU@�@0���[|�oy�T�Pf���o�G��,��y]����<N��=��i`���:�����A/.�?�0>�A���>��A��BE�8#�\�8A��<YB]��B���4��#���B�B�%��D� ia�@���zX_HEIGHYTy��M�sxB��XoA(�A�B�f@�J<��bh��ڽ@�{���w���?���A�@���@�A���q�Zpe�@?��+£�RB*�6B���B�.ߦ��l-���?An@G�1�@V���s�vT�f�� U�.0`d��hg�@���@�Y�����m?����?j��@k�{�;B��sR�@��6P@&��������,ҿ����J��(� ����;�B8)����GA�՟R� ������|iA��)���KvA9V?�	]TOOL_3�_P��}U.�j��Ż��%������r�oH�������1���������@�{��,r�,����?AZ}t
��BbRob�?�r�B��/�B���� ���Z.�A���?���Ax7��@&��o�f15����fU/�6�2����Z�Q�&��q>�u��P� �-���{�̈A�v��5����A@����@��4?<A��+_B���������B��@�j����Z������W�B���A�Z��Aa���Q�JOB_DBL_�S68�e� ������H=����<��c=F��=�����o���>ɀ�_DA��@��@É�>��h�Z���KB���� 9B��B����Q�0�����[��B,�@��mMAPF�ǥ�(﾿o/  �U0Dw�%a@���Ⱦ���?��I?a����6��������WO�AF���Y�L���@����������b@�F9��(�6�����B�C�C{8ǐi���� B
h�A�^�ATD�����L/_C?� 5�CƐ�̎F9��qW9��~��rS�d7�A�"N�����?��+^��� ���
]A
����u�BWLBu���B�Ʃ��ļ�������B�t��C��A|� ��,� ?23�oJ=Dv�%=�����:�����~>7�K��u0�P�{>�
����@=�AN�����>@J$�l@�3&=�>A��B����U�®i�B�\_�C�� �����BS�Axh=A#2���.7��v,6/i�%��!ԑ?._�<���p�~=>��>��͸��@`��i�_@���?e`�)����%����Z��A��1�.��B=�Bb��BeƠ�I��G���1��+�5A�����AZ��@����O�O�F2�%?��hz��V5���`�?��N��?B�� �4�9p���.AIڐ��Ơs@�:�@�^���p��@Ç��Z���5UB/�_�B�I[tP6z��4��)B�$y�@�OAS ���6ʜ_�����_!�hHG�;���/����:l*�)��`��!�1#A�4�	?3����@��\����@��"��]+�,�B2�ǸB�:Hm@�X��O�B�<wJ@�bAS�����po�_g�R;0F��H�<0v�=ᩋ�eP-X�=�&��)�HX
.���i�OA��5@<�� @?�d�7�=�@�q���(P����NB3B��h�D�\��i���B�@[A�=��@uB|ROS�_MOVESM_WILDER d���U6���%�y_G9����e�մ���L�W���A
�K?h�0?"��)�,4xN��A�����R�A��U�B|ӴB�?��N�X
-p���9wBA�=�A!��@�?[/��#7#�0F�1��<��!>6��y�ѺqW:~�� ��d�X
����ܕ@��\�@5�@���?������Ȕ@�o���4C�����B�pR�B����-�c��V*����aA��9@����A_�2��o"���2_DROPOFF]���7$�.b��� V5>EI��:���տ�v��:�%:����Y@���@���@��'?��zک�*@��Q�C�ό�����Ŕ���Y��\����$��A�6T@���JAt�������ҟ���=�)��P�ݾx�$��K$>����>��D��5��1�����A(��@+a��@�6Z�������+�[A����m��%�B��`B��� �X
i��D�A�՜3A"��Ad��@��ߔ������ 
U�
�^�%@3`�`�:e��l6�mq@�;L_A��n>�������@/Ê��R�Zڪ��A�� h�7 �B���]­^.��8�a� �������B�Aw��A�6���h�g쏂o_ς ����ѽ�_��J�h�3vf;�`�<D��|>��A��<|����A�V����A���5��B4���h��B�.�δ�t!\�� �������ci�Bj�"A�7��d�_AG�4�<�N�3�r�F��<��#m�;(b:�*�r;��;B��`���X
p�Alu�?���@\��G��&@�/�^�!X
�_�B��?��$2�B��65Bs6�B)�ǡ��\���l^µ��B��A�����B?��6Ϙ�*���J��P[1{ƿ�>���	����U=�`�����`X
?���A*Em��� �@�m���?�g@�� �|J��B�����B�.�B�ֻB�Pe����\������UB>����X�eB��I�������8w��o��P��:�6ڻ�@�O;�G������=�$�vy0��n�:R����7�@YN���bo@����l��{B�����B��,�B��CBיH�еp��.�¦��B?v�����B��W��<$����2��������2�H��	Fᾅ���	�=6t�)��6Β�A'@>�ۇ}@����hA����l���B����B�-��B��B�Z��вp� ����}��B1�������B�=Z�g�ˌ���2 .������;�=�P�=1����a�<�W�;�ԟ9;�TJ)@��Ҿ۴l@�T�W�ţU@�&�����B��{��B��+�B��B�O�УJ@9��WtA������j�B�N��=�62dI���
6�%<�?��@�?}�6���GS+>���@D����2���g��A_ +>	`��0����-���Z���E������B���B���A�^��Ц(*��)x��B!���U��@�q�@5d4��8ZcmL�����~�w�Y�� �K@I�h�����2w���@CzA�s��������A@y@�p����@��B��v���B��%c�8<��&����БTJ+
0���B���A���*�Y���J*SCI_�TAIL_SWI�T7U�*��Lջ�ڼ��r����oH}�@�;��S:��@�"AOX����APK_����?� ��2����aB6�?��XR!B����B�BB9�!�Ѓ�zA�V�®��B����=��B-�����l�/�)~���]U�D��VG��?Z���T��?�$�����@:o?8=�*����zv�AR��W�g%2@a�<��Em<m@��z�QtA*����)��B�0[�B���A%J��~ʅQ)�mB�(e���rD@g(��/��41�?�7(GeU:��� �@G�:��ǰ:�B��`$]�w����L�A7��f�ICm���7��٘<i����t�B9���V�B�A�B�D�B7�h���{p���y�����A�$Q�%���A}�HA��ע�FAVIZ�*��O}\T���
��;��:�P\�-0l��d�Z}�ż�@w*��I�}>I0@��Ѿ�l�����A�����2B��1�B�NB���Ǣ�R���q������A-x����4A]����8+�O"�Oo � T��n���������e�=�۫�'�޾ί��;��A�,�-�} X��o?_@�pP�� �z�p��A�M����QBDA?B��M�B�LM����Z�!hŭ�B&�2�4r\�B������P,o>o#bbo���lf��{���6�=�9���1�E���/��^�:�A�8 ���a������@�a����`�A�k������BD@�B�P�B�O��n���q�B�*y�&b�B�����C�_erhjI[m����dq��TX~�X��(��B���?�z���~����,�6�iǿ��U��4M�?��_<?b�T=����9���0��^@���]���r����Ê>����L�AVb�1p,B��XB��B�n_������R��-I�A�=k���+A��@�XZ��rw��Zhוe��~�a9���H�	�� /���A�X{غ�s�����پAW�A�P��<B?���@�i_���>�A�h�B`��Y�I��A��
�BI�B��G��̐X�Z���{�3�B/�%���AϿ!�����|��CLAMP G |m_u�T�;⤰�p"�?���d@�X@��~?03X������R��p�3J���	�`@Ml���|==��@�/�@�Z���A@Ӭ+���tB��ZB���B�C!�炻�X��p�����@�_?}�A2��N��|�RIVET�LOCv?�
7T��Nर�b�{5����"��gE���T�?U|O�?���ĽA����U�A4�	@�6Z�����Aߦ?	������A[�C�U���¦��B�f_[B�)������|����A�쭟@יCA1u�@^-b|��TOOL_2_�D���T�&W�L�@0Bþ���ܿD^�����?>���>���)�
M�����{	AY��HA��?���L?��O�������A-t�}�`=LB��{tB���Ǐ���X�B�b;���e#Ab ��wlA�}��%��;JOB_3DB�0��57χU�T�Dո��Q����`S��Qϻ��,�Q�?=ք�LSP@����?�`�@���`>�X����A�O	y��>���B��B����C�������C�A��J��[A�?Ec���P�b��x��R�䅊Q>�  �=���;��W�=�&����8=�5@�#��@�h��}�`1@� �=}�@���B@���W��c��`�BO��B���=�/�
=v�9��A���-�QA��L���q�|��qVI9S��Wk���F���=�$X<�����(<��<���:�m�������B?����=�P��Q=(�~���o�B���y��Bh���B��B����`�X�>�� ��XA��F����rA[�@�]�t�rc�Zh���5�i�t��@�-Tn��;?���@ʽ�_+�SEۚ@�p��wqHA�_���	����#x�@���@�A��
��p���d7���Y@��&�A�iwB�c�ǥ�|���"���>`���Axɖ��й�$���POS��H�Tn��T��3����]~ @�0��I��@"vo@)`����G��S��h*%��G�A�2<I�U�U�1��@���Ԯ������/T��@��BF;B�s}SB�#����V���*���+B��{'G@��51q$��6� �PV�$?SERV_M�0���H�B��Q,OU�TPU9 9��P@,RV �2X�  E (�,��PҜI�SAlQZFTOP�10 2x wd � .hbw  /��  8䀩rP�$i$s�1�%�`�  	|��6 &�P"<r  
���@ *�X�d/v/�/�/�/ �/�/�/�/??*?<? N?`?r?�?�?�?�?�? �?�?OO&O8OJO\O nO�O�O�O�O�O�O�O��K�YP�HFZ�N_CFG X�E�U�2Q?GRP 2 <W� ,B j�|POQ�D;� Bj���  B4NSR�B21�HELL�5R!X��И�SW�_�[%RSR �_�_o@o+odoOo�o so�o�o�o�o�o�o�*N_}!!fy�Q �+!���tz!gOP��r�p#�I�q�df�}�VHK 1"�[ �W�a�[��� ������͏����� >�9�K�]���������~�\OMM #�_����RFTOV_E�NB7��5�OW_REG_UI��IIMIOFWD�L��$�UJ�WAIT��TRr�Rr6�o�TIM6�7����VA6��>��_UNIT��v�LC/�TRY6�����MB_H�DDN 2%x S���LUQ�-�r� 1�m���������ٿ����2�ON_ALIAS ?e��heT�f�x� �ϜϦ�P��������� ��#�5�G�Y�k�ߏ� �߳����߂����� 1�C���g�y���H� ��������	���-�?� Q�c�u� ��������� ����);M�� q���R��� �7I[m *������/ !/3/E/�V/{/�/�/ �/\/�/�/�/??�/ A?S?e?w?�?4?�?�? �?�?�?�?O+O=OOO �?sO�O�O�O�OfO�O �O__'_�OK_]_o_ �_�_>_�_�_�_�_�_ �_#o5oGoYoo}o�o �o�o�opo�o�o 1�oUgy��H ������-�?� Q�c����������Ϗ z����)�;��_� q�����@���˟ݟ� ���%�7�I�[�m�� ������ǯٯ����� !�3�E��i�{����� J�ÿտ���϶�/��A�S�e�w�"��$S�MON_DEFP�ROG &������ �&*SYSTE�M*~���@"����RECALL �?}�� ( �})���1�C�U�g� �όߞ߰������� y�
��.�@�R�d��� ���������u�� �*�<�N�`������ ��������q�& 8J\������ ��m�"4F X�i����� �{//0/B/T/f/ ��/�/�/�/�/�/w/ ??,?>?P?b?�/�? �?�?�?�?�?s?OO (O:OLO^O�?�O�O�O �O�O�OoO __$_6_ H_Z_�O~_�_�_�_�_ �_k_�_o o2oDoVo ho�_�o�o�o�o�o�o yo
.@Rd�o ������u� �*�<�N�`������ ����̏ޏq���&� 8�J�\�������� ȟڟm����"�4�F� X��i�������į֯ �{���0�B�T�f� ����������ҿ�w� ��,�>�P�b����� �Ϫϼ�����s��� (�:�L�^��ςߔߦ� ������o� ��$�6� H�Z���~������ ��k���� �2�D�V� h�������������� y�
.@Rd���������t��$SNPX_AS�G 2&����� � 0t%|/x ?���PARAM �' ��	Ptx �3�� ���� OFT_KB_?CFG  t��OPIN_SI�M  ���/#� RVN�ORDY_DO � ��"QS�TP_DSB��a/�SR (� � & �ROS_WILD�ER LL AVE H � SS��t	� TOP_?ON_ERR*/�~�!PTN �0�A�"R?ING_PR� ,/�� VCNT_GP� 2)�x 	]/\?x J?�?n5��
�?�4�VD>10RP 1*X�p1!�?�?�?OO *OQONO`OrO�O�O�O �O�O�O�O__&_8_ J_\_n_�_�_�_�_�_ �_�_�_o"o4oFoXo jo|o�o�o�o�o�o�o �o0Bifx �������� /�,�>�P�b�t����� ����Ώ�����(� :�L�^�p��������� ʟܟ� ��$�6�H� Z���~�������Ưد ���� �G�D�V�h� z�������¿Կ�� 
��.�@�R�d�vψ� �Ϭ����������� *�<�N�`�rߙߖߨ� ����������&�8� _�\�n������2�PRG_COUN�T��2��EN�B?��M��_�UPD 1+�+T  
��t^�p� ��������������  ;6HZ�~� �����  2[Vhz��� ����
/3/./@/ R/{/v/�/�/�/�/�/ �/???*?S?N?`? r?�?�?�?�?�?�?�? O+O&O8OJOsOnO�O �O�O�O�O�O_�O_ "_K_F_X_j_�_�_�_ �_�_�_�_�_#oo0o Bokofoxo�o�o�o�o��o�o�o��_IN�FO 1,L�s2�Tp	 +�oZ�~��y� �9W�nv����D#B�Y/BX�z���VĴ�&��� �D�L�Ī-��C~�@�Q��A��B:�J�"��������/D`�A<�nA*M�9����WRE��TROL  L�1��%p��yTp����;�YSDOEBUG��M��#p�d5���SP_PA�SS��B?��L_OG -IvV��  #p��?�3װ#p(  p�qUD1:\ㄼ���_MPC� Q���!�+�27�~I�SAV .쉰���q�l�+�S�V��TEM_TI_ME 1/�W� 0 �s�]v~�
���w�s9b��MEMB/K  i���xy�����X|2�g� @��sн� �򬶯�"�3��� �{@�Y�k�}� ��ɔ����̿޿��� ��:�L�^�p�@�ϔϦϸ��ϼ�e�� ���"�4�F�X�j�|� �ߠ߲����������`�0�B�T���SKP��U���d����ﬦ	%��  v��ϯ��#p ����4�A��(5�	�'�A�`W�����tp����#p ��������2&�V�V{����#pU����! 3EWi{��� ����////A/�S/e/Y�T1SVG�UNSPDͅ '����� 2MOD�E_LIM 0�	����$2� �!1�썃%ASK_OPTION��i�a��!�_DIƀEN1��&���1BC2_GRP 22w巃��N?(#p@G C��!�G02CFG �4=;j���l��:`�?��?�?O'OO KO6OoOZO�O~O�O�O �O�O�O_�O5_ _Y_ D_i_�_z_�_�_�_�_ �_�_o1otlKo o~o�oomo�o�o�o �ozw�2o�p6 \J�n���� ���"��F�4�j� X���|���ď���֏ ���0��@�B�T��� p�[`����Ο���p� ��&�L�:�p����� b�����ܯʯ ��� �$�Z�H�~�l����� ƿ��ֿ��� ��D� 2�h�V�x�zό��ϰ� �Ϝ����.�@�R��� v�d߆߬ߚ������� ����<�*�`�N�p� r����������� &��6�\�J���n��� ������������" F��^p���0 ����0BT "xf����� ��//>/,/b/P/ �/t/�/�/�/�/�/? �/(??8?:?L?�?p? �?\�?�?�? OO�? 6O$OFOlOZO�O�O�O �O�O�O�O�O __0_ 2_D_z_h_�_�_�_�_ �_�_�_o
o@o.odo Ro�ovo�o�o�o�o�o �?0N`r�o �������� �8�&�\�J���n��� ����ڏȏ���"�� F�4�V�|�j�����ğ ���֟�����B�0� f�~�������үP� ����,��P�b�t� B����������ο� ��:�(�^�Lς�p� �ϔ϶����� ���$� �H�6�X�Z�lߢߐ� ��|������ �2�� V�D�f��z�������$TBCSG_�GRP 25����  ���� 
 @L��������/��?�  Q�c�M���q�Ы�������7��d� ���?��	� HD)̽���
>� ����cB��'4	Dp�����RG A��46K���3330���� BH|��Cj����B�B�����p:��G;�N��fff6�T�@ �������� / /��H/e/t+J(����	V3.00~t"	rc0lt#	*� �$���$�z*��  ��G  p&J) � C��(�$�?��"�#�� Ca�/9?@3��J2���8��@?L8CFG7 :������v:����"�<�<��?�?�:���? %OOIO4OmOXO�O|O �O�O�O�O�O_�O3_ _W_B_g_�_x_�_�_ �_�_�_�_oooSo >owobo�o�o�b�o �o�o�o�oE0 iT�x���� ���/��?�e��� �������ҏ ���,��P�>�`��� t�����Ο������ ��L�:�p�^����� ����ȯ�ܯ� �6� H��`�r�������� ؿƿ��� ��0�V� h�z�8ϊόϞ����� ��
��.���R�@�v� d߆߈ߚ��߾����� ��<�*�L�r�`�� ������������� 8�&�\�J���n����� ����������F 4VXj���� ���B0f Tv���z�� �//>/,/b/P/r/ t/�/�/�/�/�/?�/ (??8?^?L?�?p?�? �?�?�?�?�?�?$OO HO6OlO~O(�O�OfO dO�O�O_�O2_ _B_ D_V_�_�_�_n_�_�_ �_
o�_.o@oRodoo �ovo�o�o�o�o�o �o*N<^`r �������� $�J�8�n�\������� ��Əȏڏ��O(�:� L���|�j�������֟ ğ����0�B�T�� x�f�������ү��� ��¯,��P�>�t�b� ������ο����� �:�(�J�L�^ϔς� �Ϧ����� ����6� $�Z�H�~�lߢߴ�^� ����d��� ��D�2� h�V�x��������� ����
�@�.�d�v� ����T����������� <*`N�r ������& 68J�n�� �����"//F/ ����p/�/,/Z/�/�/ �/�/?�/0??T?f? x?�?H?�?�?�?�?�? OO,O>O�?bOPO�O tO�O�O�O�O�O_�O (__L_:_p_^_�_�_ �_�_�_�_�_o o"o $o6oloZo�o~o�o�o �o�o�/&�oV Dzh����� �
��.��R�@�v�8d�����  ��ă� Ć؏Ă�$�TBJOP_GR�P 2;����  ?�/  C4Ă	�����=��䔀L���X���Ą9�&X�^,^XĄ @�����ߐD)�t�CQ?p�D5mą�x��i���>�����ަ�<ѥ�t�?3�33?W
=̑Bp  A�����yDِ�C���xj�͑͐>���$��6�<�~��?L�B�uԒ�  cBޟ��K���CQff�6������Ǫ<������ಐ]�h�	�ąCj�9�$����S�����A�S�;���B�̚ݐؑ�����$�6�Ȧ]�տ�<�ex�fff?�+=q����� ��/��;�ND���S�͑<e�w�<?�x������C�������ϐ� ������������K� &���j߄�n�|ߪ��� ��p�������:�k�����Ć�  0���	V3.00��rc0lI�a*��I���ĄB�r��  F�� �F�P F�� �F�` G � �G� Gp �G@ G'� �G/� G;� �GG8 GO �GZ� Gb� �GnH Gv �G����� G������F�F�F�z  F�� F�� F������� F�  G�.���� (�7�� G?h GK�  =aG�=#��
T�h��� ��Ώ����Ć��?�A�h�<��ESTP�ARW���	��H�R ABLE 1�>�� ��ăD���� 8p��������Çˁ��	��
�����Yā�������6RDIA�Xj|���O"4>PbHt�:S � �
 G/Y/k/}/�/�/�/�/ �/�/�/??1?C?U? g?y?�?�?� #/� W�9����������:�2NUoM  ���d�̀ V :_CFG ?�K�ZCh�@��IMEBF_TT%UE�����FVER�1V��CR 1@I �8��PY��bQ ���?  J_\_n_�_ �_�_�_�_�_�_�_o "o4oFoXojo|o�o�o �o�o�o�o0�B~��3ZlHz�xq���B~{�<���B~UTU�!�_�DE6�H�B~OTF8n���B~$C����B~$W���H{C8�,�HzRIDN�`�R/T_�AV@&U MI_CHAN�G� &U ɓDBGL�VL�G&U̐E�THERAD ?�)����0�(�:e+�4:55:bb:26 (�m7;�28O�29�oROUTP!��!~���	̐SN�MASK�&S%�255.ڥ��د������ OOLO_FS_DIW������ORQCTRL� A9[���z�T i�����¿Կ���
� �.�@�R�d�vψϚ� �Ͼ���h������;PEk�TAI�?��PGL_CONF�IG G�I�A���/cell/�$CID$/grp1ߏߡ߳�������C��&�8�J� \��߀�������� i����"�4�F�X��� �������������w� 0BTf��� �����s�@,>Pbt�>}	 �����/rA�,/-�a/s/�/�/ �/�/�/�/??'? 9?�/]?o?�?�?�?�? �?X?�?�?O#O5OGO �?kO}O�O�O�O�OTO �O�O__1_C_U_�O y_�_�_�_�_�_b_�_ 	oo-o?oQo�_uo�o �o�o�o�o�opo );M_�o��� ���l��%�7��I�[�m�hдU�ser View� }�}}1234?567890���� ԏ��� ���]� �����2���b�t�����������-���3 E�
��.�@�R�d�ß��3�4����Я��� ��w�9�3�5��r� ��������̿+��3�6a�&�8�J�\�nπ�߿��3�7�������@�"�4ߓ�U�3�8�� �ߠ߲�������G�	��� lCamera����N�@`�r����EA� ������"�4�F�X�j�`�  (�D�=� ����������8 J\����������(���q&8 J\n�'��� ��/"/4/F/� �����/�/�/�/�/ �/�?"?4?/X?j? |?�?�?�?Y/���K?  OO$O6OHOZO?~O �O�O�?�O�O�O�O_  _�?)�ɵOj_|_�_ �_�_�_kO�_�_oW_ 0oBoTofoxo�o1_� ��!o�o�o�o0 �_Tfx�o��� ����o�|ٍB� T�f�x�����C��ҏ �/���,�>�P�b�	��9���ǟٟ ������3�E��V��{�������ïկd�	*�0[��"�4�F�X� j��������Y�ֿ� ����0�ׯ�/�1� Կ�ϛϭϿ����ϊ� ��+�v�O�a�s߅� �ߩ�P�*��@���� �+�=�O���s��� �߻����������� ��	��a�s������� ��b�����N�'9 K]o�(�:�u+ ���'��K ]o������ ��:��;�9/K/]/ o/�/�/:�/�/�/&/ �/?#?5?G?Y? /:� M[�/�?�?�?�?�?�? �/#O5OGO�?kO}O�O�O�O�Ol=   p9�O__*_<_N_`_�r_�_�_�_�[   }�I?��B�  �Q�]�Y�_o$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh z������� 
��.�@�R�d�v��� ������Џ�����*��^  
l0( � ��@( 	 <�r�`��������� ޟ̟���8�&�\��J���F��Z � Oůׯ�\O��1� C�U�g�n3�������� ��ٿ����!�3�z� W�i�{�¿�ϱ����� ����@��/�A߈�e� w߉ߛ߭߿����� ��`�=�O�a�s�� ���߻�����&��� '�9�K�]�������� ����������#j� |�Yk}����� ���B1C� gy����� �	/P-/?/Q/c/u/ �/���/�/�/(/? ?)?;?M?_?�/�?�? �?�/�?�?�?OO%O l?IO[OmO�?�O�O�O �O�O�O2ODO!_3_E_ �Oi_{_�_�_�_�_
_ �_�_oR_/oAoSoeo wo�o�_�o�o�oo�o�+=O�ov�@� qr~��qs�xw\���)frh�:\tpgl\r�obots\r2�000ic�u_210l.xml^ ��*�<�N�`�r�������������ُ� ���!�3�E�W�i�{� ��������՟���� �/�A�S�e�w����� ����ѯ�����+� =�O�a�s��������� Ϳ߿���'�9�K� ]�oρϓϪ������� �����#�5�G�Y�k� }ߏߦϠ��������� ��1�C�U�g�y�� �ߜ���������	�� -�?�Q�c�u������x��a x�p<�< �p ?� ����������$
, Z@r�v��� ���&D*<�^��f�`(�$�TPGL_OUT?PUT J�a�aw� � ��//)/;/M/_/ q/�/�/�/�/�/�/�/ ??%?7?I?[?m??������2345?678901�?�? �?�?�?�?C�b�?-O ?OQOcOuO�OO�O�O �O�O�O_�J}_7_ I_[_m___)_�_�_ �_�_�_o�_oEoWo io{o�o%o�o�o�o�o �o�o�oASew ��3����� ��'�O�a�s����� /�A�͏ߏ���'� ��5�]�o�������=� ��۟����#���͟ Y�k�}�������K��� �����1�ɯ?�g��y�������G�� $${�?��� �	�;�-�_�Qσ�u� �ϙ��Ͻ������� 7�)�[�M��qߣߕ� �߹������}��)�@;�M�_�q���@��������� ( 	 �����#��G� 5�k�Y�{�}������� ������1Ag U�y��������-Q�6� ? <<� ��u����/ �:r8/J/�V/�/Z/ l/�/�/&/�/�/�/�/ 4?F? ?j?|?�/d?�? L?�?�?�?�?O0O�? OfOxOO�O�O�O�O �OBOTO_,_�O4_b_ <_N_�_�__�_�_z_ �_o�_oLo^o�_fo �o.o�o�o�o�o  po�oHZ�o~�j ��$����2� D��0�z����� \�Ώ��ҏ�.�@��� D�v��b�������� ��R�ܟ*�ğ�`�r� L��������ޯ𯊯 �&� �2�\���̯�� ��>���ڿ��ƿ�"� ��F�X��Dώ�h�z������h)WGL�1.XML�����$TPOFF_L�IM m��i���N_SV�!�  ��3�P_MON KeS5ԣ���2��STRTCHK �Le3�&��VTCOMPATH����7�VWVAR �Mh���L� ��� ��{���_DEFPRO�G %��%
�ROS_WILD7ER _�H l���_DISPLAY�(З�=�INST_�MSK  �� =y�INUSc����<�LCK���QU?ICKMEN���oSCRE�e~��t_sc�`��/�4�3�E�ST���3�RACE_CF�G Nh����}�	�
?���HNL 2OL�E���� "�����0�BTfx
��ITE�M 2P�� ��%$123456�7890��  �=<���  #!��X �y���� 7I/m-/�=/c/ ����/!/�/E/ �/?)?�/M?�/�/�/ O?�/�?�?�?A?�?e? w?�?O[O�?O�O�? �OO+O�OOO_sO3_ E_�O[_�O_�__�_ '_�_�_oo_o�_�_ �_1o�_�o�o�o#o�o GoYoko�o�oas �o�o�1�U �'��=������ ��	���ۏa�Q�c�u� �������i������ ş)�;�M�ǟq��C� U���a�ݟ����ӯ 7���	�m������l� ǯ��믫���!�ӿE� �� �{�;ϟ�K�qσ� 翏���/ϩ�S��� %�7ߛ�[߿�����g� ������O���s߅� N��i��ߍ����P'�9����S��Q��>��  ��� ��^�U�
 �k���x���6�UD�1:\�����R_GRP 1R��� 	 @ ^�	?-cQ�u�� ��
������
�?�   %7!WE{i� ������//�A///e/S/u/�/	���/�/�SCB ;2S#� ? ?1?C?U?g?y?�?�?��UTORIAL� T#����?�V�_CONFIG sU#��� %@���?MO�7OUTP�UT V#�8@��SO�O�O�O�O �O�O__'_9_K_]_�o_5A�\Reg�ular Opt�ion\R632� : KAREL t_�_�_�_�_�_o!o 3oEoWoioU�ЄO�o �o�o�o�o�o) ;M_q�T�o�� ������,�>� P�b�t��������Ώ �����(�:�L�^� p���������ʟܟ�  ��$�6�H�Z�l�}� ������Ưد����  �2�D�V�h�z����� ��¿Կ���
��.� @�R�d�vχ��ϬϾ� ��������*�<�N� `�r߃ϕϨߺ����� ����&�8�J�\�n� ��4E/�(O�O������ ��
��.�@�R�d�v� �����߾������� *<N`r�� ������& 8J\n���� ����/"/4/F/ X/j/|/�/�/��/�/ �/�/??0?B?T?f? x?�?�?�/�?�?�?�? OO,O>OPObOtO�O �O�O�?�O�O�O__ (_:_L_^_p_�_�_�_ �O�_�_�_ oo$o6o HoZolo~o�o�o�_�o �o�o�o 2DV hz����o�� �
��.�@�R�d�v��������������̏ޏȁ��	����\Regular� Option\�R632 : K�AREL ock?et Msg�]� o���������ɟ۟� ����p%�7�I�\�n� ��������ȯگ��� ��4�F�X�j�|��� ����Ŀֿ����� 0�B�T�f�xϊϜϮ� ����������+�>� P�b�t߆ߘߪ߼��� ������'�:�L�^� p�����������  ��#�6�H�Z�l�~� �������������� �1�DVhz�� �����
- @Rdv���� ���//)</N/ `/r/�/�/�/�/�/�/��/??&>�$TX�_SCREEN �1W��Ȁ�}�&?j?|?�?�?�?�?X?�W?O O(O:OLO^O�?�?�O �O�O�O�O�OeO_�O 6_H_Z_l_~_�__�_ +_�_�_�_o o2o�_ �_hozo�o�o�o�o9o �o]o
.@Rd �o��o����� �}�<�N�`�r��� �����1�ޏ�����&�8���\��$UA�LRM_MSG k?F9�S0 T� )*����џğ���� ��<�B�s�f��������o�SEV  �}��m�ECFoG YF5P1�  )%@�  }A�   B�0"�R1����@�?��R�*�4�S��B�=�U62D F5h�z�������¿Կ����
�J1��GRPw 2Z� 0<��  	 ����?Nā�p��?��7?���"?MĴ��'g�I_BBL_NOTE [��T��l�0"K02!�o�DE�FPROy�%}�� (%DATA�MAP OSIT�ION_��_��R�AM)'%TOO�L_4_PICK�_A��ACH�� %��&��J�5�n�Y߀��}߶��߳���j�FwKEY�� 1\F9�F�p �)& ��N�`�7���m�,(����)$��O?INT  ]����? ANCEL��&����NDIRECT�'�)� EXT S�TEPS�V�OUC�HUo�����RE INFO�������� ��!EW>{b�������� ��  frh�/gui/whi�tehome.pngJ\n��>!point5�����/�FRH�/FCGTP/wzcancel��O/a/s/�/�/�indirec��/�/��/??#/5 nex��/T?f?x?�?�?�t?ouchupD?�?��?�?O O+?� fo �?[OmOO�O�O�7�O �O�O�O__+_�OO_ a_s_�_�_�_8_�_�_ �_oo'o�_Ko]ooo �o�o�o�oFo�o�o�o #5�oYk}� ��B����� 1�C�_�q������� ��ˏ����%�7� I�؏m��������ǟ V�����!�3�E�W� �{�������ïկd� ����/�A�S��w� ��������ѿ�r�� �+�=�O�a��ϗ� �ϻ�����n���'� 9�K�]�o��ϓߥ߷� ������|��#�5�G� Y�k��ߏ������� ������1�C�U�g��y���� �����������,�6� INS�T ]?A IR�ECTk�% ND����CHOIC�EZ�  EDCMD�%>%b I������ �/�:/L/3/p/O���%whitehomeJO�/�/�/�/�/�<insC?4?F?X?�j?|??�0direc#3'?�?�?�?�?O <�84OFOXOjO|O�O>8choic�#3O��O�O�O�O_:edcmd0B2OK_]_o_��_�_;arwrg /O�_�_�_ oo	�6o HoZolo~o�oo�o�o �o�o�o �oDV hz��-��� �
���@�R�d�v� ������;�Џ��� �*���N�`�r����� ��/E�ޟ���&� 8�?�\�n��������� E�گ����"�4�F� կj�|�������ĿS� �����0�B�ѿf� xϊϜϮ�����a��� ��,�>�P���t߆� �ߪ߼���]����� (�:�L�^��߂��� ������k� ��$�6� H�Z���~��������� ����y� 2DV h��������ڽ���� ���/AcuO,a/�Y/�� � /�$//H/Z/A/ ~/e/�/�/�/�/�/�/ ?�/2??V?=?z?�? s?�?�?�?�?ş
OO .O@OROdOs�O�O�O �O�O�O�O�O_*_<_ N_`_r__�_�_�_�_ �_�__o&o8oJo\o no�oo�o�o�o�o�o �o�o"4FXj| ������� �0�B�T�f�x���� ����ҏ������,� >�P�b�t�����'��� Ο�������:�L� ^�p�����#���ʯܯ � ��$��?H�Z�l� ~�������ƿؿ��� � �2���V�h�zό� �ϰ�?�������
�� .߽�R�d�v߈ߚ߬� ��M�������*�<� ��`�r�����I� ������&�8�J��� n�����������W��� ��"4F��j| �����e� 0BT�x�� ���a�//,/�>/P/b/9�d+�>9�����/�/ �-�/�/�/�&,�?? �?:?!?^?p?W?�?{? �?�?�?�?�?O$OO HO/OlO~OeO�O�O�O �O�O�O�O __D_V_ 5�z_�_�_�_�_�_� �_
oo.o@oRodo�_ �o�o�o�o�o�oqo *<N`�o�� ������&� 8�J�\�n�������� ȏڏ�{��"�4�F� X�j�|������ğ֟ ������0�B�T�f� x��������ү��� ���,�>�P�b�t��� �����ο��ϓ� (�:�L�^�pςϔ�k_ �������� ���6� H�Z�l�~ߐߢ�1��� ������� ��D�V� h�z���-������� ��
��.���R�d�v� ������;������� *��N`r�� ��I��& 8�\n���� E���/"/4/F/ �j/|/�/�/�/�/S/ �/�/??0?B?�/f?�x?�?�?�?�?�?����;�������?O!M�?COUO/F,A_�O9_�O�O�O�O �O_�O(_:_!_^_E_ �_�_{_�_�_�_�_�_ o�_6ooZoloSo�o wo�o�o���o�o  2DS?hz��� ��c�
��.�@� R��v���������Џ _����*�<�N�`� �������̟ޟm� ��&�8�J�\�럀� ������ȯگ�{�� "�4�F�X�j������� ��Ŀֿ�w���0� B�T�f�x�ϜϮ��� �����υ��,�>�P� b�t�ߘߪ߼����� ����o(�:�L�^�p� ��ߦ�������� � ���6�H�Z�l�~��� ������������� 2DVhz��- ����
�@ Rdv��)�� ��//*/�N/`/ r/�/�/�/7/�/�/�/ ??&?�/J?\?n?�? �?�?�?E?�?�?�?O "O4O�?XOjO|O�O�O �OAO�O�O�O__0_�B_�D[�����m__�]i_�_�_�V,�o�_�oo o>oPo7oto[o�o�o �o�o�o�o�o( L^E�i��� �� ��$�6��Z� l�~��������O؏� ��� �2�D�ӏh�z� ������Q����
� �.�@�ϟd�v����� ����Я_�����*� <�N�ݯr��������� ̿[����&�8�J� \�뿀ϒϤ϶����� i����"�4�F�X��� |ߎߠ߲�������w� ��0�B�T�f��ߊ� ���������s��� ,�>�P�b�t�K����� ����������(: L^p���� �� �$6HZ l~����� �/�2/D/V/h/z/ �//�/�/�/�/�/
? �/.?@?R?d?v?�?�? )?�?�?�?�?OO�? <ONO`OrO�O�O%O�O �O�O�O__&_�OJ_ \_n_�_�_�_3_�_�_ �_�_o"o�_FoXojo�|o�o�o�o���k}�������o@�o}�o#5v,!� f��q���� ����>�%�b�t� [������Ώ���ُ ���:�L�3�p�W��� ����ʟܟ� ��$� 3oH�Z�l�~������� C�د���� �2��� V�h�z�������?�Կ ���
��.�@�Ͽd� vψϚϬϾ�M����� ��*�<���`�r߄� �ߨߺ���[����� &�8�J���n���� ����W������"�4� F�X���|��������� ��e���0BT ��x������ ��,>Pbi �������� /(/:/L/^/p/��/ �/�/�/�/�/}/?$? 6?H?Z?l?~??�?�? �?�?�?�?�? O2ODO VOhOzO	O�O�O�O�O �O�O
_�O._@_R_d_ v_�__�_�_�_�_�_ o�_*o<oNo`oro�o �o%o�o�o�o�o �o8J\n��! ������"�� �$��� ���M�_�q�I������,��֏������ 0��T�;�x���q��� ��ҟ�˟��,�>� %�b�I���m������� �ǯ���:�L�^� p��������ʿܿ�  ��$ϳ�H�Z�l�~� �Ϣ�1����������  ߯�D�V�h�zߌߞ� ��?�������
��.� ��R�d�v����;� ��������*�<��� `�r���������I��� ��&8��\n �����W�� "4F�j|� ���S��// 0/B/T/+�x/�/�/�/ �/�/��/??,?>? P?b?�/�?�?�?�?�? �?o?OO(O:OLO^O �?�O�O�O�O�O�O�O }O_$_6_H_Z_l_�O �_�_�_�_�_�_y_o  o2oDoVohozo	o�o �o�o�o�o�o�o. @Rdv��� �����*�<�N� `�r��������̏ޏ �����&�8�J�\�n�h����i ���i �����ϟ������,�F��� j�Q�������į��� �����B�T�;�x� _�������ҿ����ݿ �,��P�7�tφ�e/ �ϼ���������(� :�L�^�p߂ߔ�#߸� ������ ���6�H� Z�l�~�������� ����� ���D�V�h� z�����-��������� 
��@Rdv� ��;��� *�N`r��� 7���//&/8/ �\/n/�/�/�/�/E/ �/�/�/?"?4?�/X? j?|?�?�?�?�?���? �?OO0OBOI?fOxO �O�O�O�O�OaO�O_ _,_>_P_�Ot_�_�_ �_�_�_]_�_oo(o :oLo^o�_�o�o�o�o �o�oko $6H Z�o~����� �y� �2�D�V�h� �������ԏ�u� 
��.�@�R�d�v�� ������П������ *�<�N�`�r������ຯ̯ޯ���$U�I_INUSER  ���#���  ���_MENH�IST 1]#��  (�2��0)/SOF�TPART/GE�NLINK?cu�rrent=me�nupage,1�631,1 RT/_POS��1B����ӿ忋�(|���95�5����AFE_9�3��4�F�X�jό�'l ώ�74��MP���ERROR_MO�VE_PROGRAM2�����uχϑ�37��5 �Ŷ�Kߘ]�o߉�� 	��62G�TY_��G���P��}ߏߑ�5��I�� ��]�o����Ϣ����ITION_MA ��L���������;𣰾�P�b�t��� ����w�������� ���� �(:L ^p��#��� � �6HZl ~������ / /�D/V/h/z/�/ �/-/�/�/�/�/
?? �/@?R?d?v?�?�?�? ���?�?�?OO*O-? �?`OrO�O�O�O�OIO �O�O__&_8_�O\_ n_�_�_�_�_E_W_�_ �_o"o4oFo�_jo|o �o�o�o�oSo�o�o 0B�o�ox�� ����?���,� >�P�b�e�������� Ώ��o���(�:�L� ^�폂�������ʟܟ �}��$�6�H�Z�l� ��������Ưد�y� � �2�D�V�h�z�	� ����¿Կ����� .�@�R�d�vψϋ��� ��������ߕ�*�<� N�`�r߄�ߨߺ��� �������8�J�\� n���!�������� �����4�F�X�j�|� ����/����������	��$UI_P�ANEDATA �1_���L�  	��}c/frh/c�gtp/flex�dev.stm?�_width=0�&_height�=10| m ice�=TP&_lin�es=15&_c�olumns=4�| font=24�&_page=w�holem (�)�prim��  }�-?Qcu )w���� ���/ /=/O/6/�s/Z/�/�/�/�/�ߐ� �  �$ 0fr�s/optntrKeep q�2��30�1�dou�bm 2�/�(ualk?�?�$bi6�?�? �?�?Om?*O<O#O`O GO�O�O}O�O�O�O�O �O_�O8_J_1_n_�'� �#  ��ArL�9i?�3�(� A?�t�P3w_R[hirdo5oYo ko}o�o�o�oZ_�o�o �o�o1U<g �r�����	�|^,�NIoN�`�r� �������̏?o��� �&�8�J���n���g� ����ȟڟ�����"� 	�F�X�?�|�c����� %�7������0�B� ��f�ُ��������ҿ ���]���>�%�b� t�[Ϙ�ϼ��ϵ��� ���(��L߿�ѯ�� �ߦ߸�����/� �� ��6�H�Z�l�~���� ������������2� D�+�h�O��������� ����Y�k�)�.@R dv������� �*�N`G �k�����/ �&/8//\/C/�/�/ �/�/�/�/?"? u/F?�j?|?�?�?�? �?�?=?�?�?OOBO TO;OxO_O�O�O�O�O��O�O_�O,_�/�*��7_p_�_�_�_�_�_) ^_�_b5�_o-o?oQo couo�_�o�o�o�o�o �o�o�o;M4q X����[8�#�+��$UI_POSTYPE  �%�� 	 �AV�[6�rQUI�CKMEN  ���i�;�RESTORE 1`�%�%����d2������d2m ӏ��� �2�D��h� z�������S�ԟ��� 
��Ǐ)�;�M����� ������Яs����� *�<�N��r������� ��e�ǿٿ�]�&�8� J�\�n�ϒϤ϶��� ��}����"�4�F�� ��e�w��ϛ������� ����0�B�T�f�x� ������������ ����P�b�t����� ;������������:L^p�<�SC�REL�?Q��u1sc��uU2�3�4�5��6�7�8��T;AT�� ��%�zUSER� ��Sks�P3P4PU5P6P7P8P��pNDO_CFG� a�#��pP�D :��None?�1_I�NFO 2b�%�^�0%��[8 �.//R/d/G/�/�/ }/�/�/�/�/�/?*?�?N?5��OFFS�ET e�� [?#��+�?�?�?�? O�?O8O/OAO�?EO �O�O�O�O�O�O�O�O�__cKa�e]S_�_
�x_�_��WOR/K f�f_�_��_�_]?0UFRAME  ����RTOL_ABRqTLo�dbENBmo~^hGRP 1g���]�Cz  A� �c�a��o�o�o�o	 -?{`fK�U�h�~|kMSK  ����%�`fNIa%���%RIVE�TLOCATIO�N/of8R_EVN�l`�t��v�2h�};
 h�U�EVl`!td:�\event_u�ser\�0�C7�5��_% F�])�SP�.�3�spotw�elde�!C6 ��k�}�� 5T!5_D� �7�⇞q��&��j� ��J�\�՟�������� ȟA��e��"�X��� ��ѯ|���į��=� ���s������T�f�@߿��Ϯ����W�P32i;�Q8��g�y� UϞϰϋ����� ��
����@�R�-�v� ��c߬߾ߙ���������*��;�`�r��$�VALD_CPC� 2j}; 8N�� 2_��oo���,�qx#	�dS�P�Mqg�O� x������������ $6E�W�i�{�} ���������  2ASew��� ����/./� Oas�@/��/� ��//�/*?<?K/]/ o/�/�/�/�?E?�/�/ O?&O8OG?Y?k?}? �?�O�?�O�?�?�OO _4_F_UOgOyO�O�_ �O�_�O�O�Oo_0o BoQ_c_u_�_�_�o�_ �o�_�_o,>P _oqo�o)��o��o �o�%:�L�[m �����܏�� �!�6�H�Z�i�{��� ����Ï؟���/� � �D�V�e�w������� ���������+�@� R��s�������d�ͯ �����'��N�`� o���������ɿ��i� ���&�5�J�\�k�}� �ϡϳ���������� ��1�2�X�j�yߋߝ� �߱�������	��0� ?�T�f�u����� ��������,;�P bt������M��� �%:I^p ������ / !6/EZ/l/~/� ����/��/// S/D?3?h?z?�/�/�/ �/�/�/�?
O?+?@O O?dOvOO�?�?�?�? �O�?_O'O�OKO=_ r_�_�O�O�O�O�O�O o�_#_5_JoY_no�o �_�_�_�_�_�o�_ o1oUoV|��o �o�o�o��o�- ?T�cx������ ������)�;�P� _�t���������ˏq� ߟ��%�7�I�^�m� ��������ǟٟ� � �$�3�E�Z�i�~��� ����ïկ��� � /�A�w�h�WόϞϭ� ��ѿ����	�.�=� O�d�sψߚ�1߻��� ���Ϭ��*�9�K�� o�a��������������$VARS�_CONFIG �kL�3��  FP����CCRG_C_FG n3�% ���D���B�H  Ap����Ce��������?���z���=������A V�MR_GR�P 2t3�����	��?�  %�1: SC13?0EF2 *?C ���L�������e5�����A@��;CȌ� 	������&�)�A���F����f� B��́�� ������/� 6/!/3/l/�M/�/�/��/�/��/?T�TC�C_�u3�����@9E��#�G�F(�a�2v3��s�234567�8901}?�2��3���%�M�?�8�����!3��?�7B��0�������:�o=L� ��|,@|?�����}���nM0As��O�?�3 �O�O�?�?�?O"O4O FOXOjO|O�O�_�O�O �_�O�O o_0_B_T_ }ox_�_�_�o�o�_�o o*o@>oPoboto��o�o�o�c\4MOD�E  ?�;� �\4RSLT w3���%"�?�?A��/ J�w��k�3���a\4?SELECT�s����yIA_WOR�K x3���<]���,		M�B>%�G�P �<�<���SIONTMO�UԄ!r;��  ��O�_�y������l;1 �FR:\Q�\DA�TA\�� ��� MC��LOG���   UD1搖EX���' B@ ����Ց  Pendant�̚&�J������� n6  ��������-�|s���   ���䙠֐��TRAcIN��� 
��3p�����������@�L�p�z3� (�!�<��)<�F� X�j�|�����ֿĿ޿������0��ISSTA�{39,� �ϡϳ��$����m��_GE_�|3��`��
]�[���H�OMINb�}�?������rq�rq��C�7�����J�MPERR 2~3�
  �o�� u5����������� !�3�E�[�i����X3����REb�|ή�LEX Ԁ��1-e��VMPH?ASE  ��s��r��OFFSE�T_ENB  ^�$VP2w��@Х0@МDӡ���@�F����'p?s33�������T͔��P��v|$1�Є���٣�m� E����[1�����_�3���A7���ڤs�\�i�!�A�'�4P����3����Cܪ5�>� �������f�� H=a�} �l~ ���J�"/)/ XJ/�V/�/z/��/ ��//?0/B/�/2? @?R?h?�/�?�/�/�/ �??�?v?O*O<OfO �?�?hO�?�O�OO�O `O_,_&_pOe_�O�_ �O�_�O�O8_�_�_�_ oZ_Oo~_�_�_�o�_ lo"o�o�o�oDo�o zoo��o�� ���@2�dY� �����������·���TD_FILTuE�Ѕ� ԰�����i�0�B�T�f� x���������ҟ��� ���#�5�G�Y�k�}��������SHIFTMENU 1���<��%������ݯ �<��%�r�I�[��� ������ǿٿ&�����\�3�	LIV�E/SNAPP�?vsfliv�n�����ION �S�U����menu �Ϭ�F���ׂ��t�����MOt���z��ZD<ԉ����< �`��$WAITDIN?END  +�@��Pҥ�OKZ���OU�T����S����TI]M����G�� <���_���?��?�,���RELE2�[��سTM��L����_GACT��Z�8��w�!�DATA ���9�%ROS_�MOVESM_WGILD��p�H�!��RDIS�����$XS>ҋ�٤�t����  ��XVR�>��f��$ZA�BC_GRP 1]��� ,L�2v����~�(�VSPT ��f���H�

�
߀�ʍ�B_DCSCH@ЏP�pb��	��ZIP=����N�?Qc�<
MPCF_G ;1��� 0u�M�ȳy�v�p�u�� 	�������  ?�-��?8 ���u�5[?�1Ҋ>��>�GX'<hN!?�{yD�L���-�C~�H�����:B����#����?���d?q�齫?G�Ĵ�&/$&�n.'�: &<hKM�B,�R/d"cj/�|(��//�)?!�� �������/D`�A�<oA*P��9�F<�V0sZ0I^2?8�0�?�?�?�?@�?�;~/�/�/�"��/��/��@ГWD_�CYLINm�2��� �!� ,(  *�O�M(��O0�O�O_�M  ?=_ O_a^�O�_�O�_�_�_ �_!_oo&oi_Jo�_ �_�ogo�o�o�_�o�o�;�2�dG;�w�� �7l�?m?��|h'�!���qA�wD�SPHERE 2��M�>o��o�P� 7�t��o�����8o�� �e����:�!���p� ��ɏۏ��+�ܟß՟��Y�6�H�Z���ZZ�� �L�