��   >D�A��*SYST�EM*��V9.3�0146 5/�27/2021 A 
  ����CELLSE�T_T  � w$GI_ST�YSEL_P �7T  
7ISO:iRibDiTRA�R|��I_INI; �����bU9A�RTaRSRPNSS1Q23U4567y8Q
TROBQ?ACKSNO� �)�7�E� S�a�o�z�2 3 4 5* 6 7 8aw.n&GINm'D�&� �)%��)4%��)P%���)l%SN�{(O�U��!7� OPT�NA�73�73.:BP<;}a6.:C<;CK;�CaI_DECS�NA�3R�3�TR�Y1��4��4�PTHCN�8D�D>�INCYC@HG��KD�TASKOK�{D�{D�7:�E �U:�Ch6�E�J�6�C�6U�J�6O�;0U��:IATL0RHaRbH<aRBGSOLA�6�VbG�S�MAx��Vp��Tb@SEGq��T��T�@REQ �d�drG�:Mf�G�JO_HFAUL��Xd�dvgALE@� �g�c�g�cvgE� x�H�dvgNDBR�H<�dgRGAB�Xt�b���CLMLI�y@   �$TYPESIN�DEXS�$$C�LASS  ����lq�����apVERSION�ix  �1b�$'61�r���p��q�t+ �UP0 �x�Style Se�lect 	  ���r�uReq. _/Echo���y�Ack�s�sI?nitiat�p�r��s�t@�O�a�dp���	��  ��U��������:q�������q��s�Option b�it A��p�B�����C�Deci�s�cod;��zTryout mL���Path se}gJ�ntin.��II�yc:��Ta�sk OK��!�M�anual op�t.r�pAԖB�ޟԖC�� dec�sn ِ�Rob�ot inter�lo�"�>� isSol3��C��i/�<"�z�ment���z�ِ����_�sta�tus�	MH ?Fault:��ߧAler��%��pn@r 1�z L���[�m�+�; LE_�COMNT ?>�y� � ��� ��Ŀֿ�����0� B�T�g�xϊϜϮ��� ��������,�>�P�@b�t߆ߘߪ߼��� ��������)�;�M�_�q�������4t������ch�� ���/�A�S�e�w���ܮ����4�� ���������� w �;���bL� $M#q���TM_�����߽�� mp��7I [m����� ����
B/T/f/x/ �/�/�/�/�/�/�/? ?,?>?P?b?t?�?�? �?�?�?�?�?OO(O :OLO^OpO�O�O�O�O �O�O�O __$_6_H_ Z_l_~_�_�_�_�_�_ �_�_�$//0oBoTo go�o�o�o�o�o�o�o �o@>/$o:L �������� �(�:�L�^�p����� ����ʏ܏� ��$� 7�\�Z�l�~������� Ɵ؟��� �2�D� V�h�z�����į¯ԯ����
�j��U�� ���  Ȑ�E�NAB  ����������ȿڿ� ���"�4�F�X�j�|� �Ϡϲ���������߀�0�B�T�f�xߊ� �СҎ߸�������  ��$�6�H�Z�l�~�x���Q�MENU^��i���NAME {?%��(%$*���?�o{%	NORM?ALIZE ����_TO_VI�S%��L�ION� ���L�H�DR�ILLO��CL�AMP ���U�N������_HEIGHT��>�Y��PON���RI�VETLOCAT�o�F��:H��T�OOL_2_PI�CK_APROA�CH � ��	L�EAVE ����DROPOFF�������3@��N�6�3��3USAFE�_POSIeO
T�RANSPORT`��S���TY!/�SD�:�
MANGTEC/<� 1R �/��$��1��:�/�	4�/�/V7��4
??�:;?�p��000�  %�JOB_DBL�_�1OfpSETrL2-OfpARML)3UOdrUL4Ofp��4AM5�OfpXS�EL6�OfpORGrL7�Ofp�4L�8_csL9H_TT KO|_&A)O�_&AQO �_&AyO�_&A�Oo&A �ODo&A�Olo&A_�o &AA_�o&Ai_�oNA�_ NA�_4NA�_\NA 
o�NA2o�NAZo� NA�o�NA�o$�NA�o L�NA�ot�vA"��vA31 ��Ə_3r�vA3ۏ�w@�<�vA �d�vA���vA:��� vAb�ܟvA����A,� ,��AJT��A�|��A ����AR�̯�Az��� �A����AʟD��A� l��A����AB����A j���A����A��4� �A�\��A
����A2� ���AZ����A�����A ��$��AҿL��A��t� �A"Ϝ��AJ����Ar� ���A����A��<��A ��d��Aߌ��A:ߴ� Qb���Q���Q�� ,�Q��T�Q�|�Q *��QR���Qz��� Q��Q��D>Q�� l>Q��>QB��>Q j��>Q��>Q��4 >Q��\>Q
�>Q2 �>QZ�fQ��fQ �$/fQ�L/fQ�t/@fQ"�/fQJTTļ�O�/�":/VRUF�_RIVETLO�CA�2T?WQD1E�GENFRAME R?<5T�?�?_�,?�USCOGNEX�_ERROR_M�OVE_PROG�u0M[NORMA�LITY�?�8%*4D�?NZ3OlOWO�O�{O�OOY
ROS_?WILDER�O�O �O�O�O7_"_[_F__ j_�_�_�_�_�_�_�_ !ooEo0oB`�OWoAo {o�o�o�o�o�o�o /AS�w� ������.�� R�=�v�a�s������� ���ߏ��<�'�9� K�]���������ޟɟ ۟����#�\�G��� k���������ů��� "��F�1�C�U�g�y� ��Ŀ���ӿ���	� �-�f�Qϊ�uϮϙ� �Ͻ�������,��P� ;�t�_�q߃ߕ��߹� ��]n�<$�