��   8��A��*SYST�EM*��V9.3�0146 5/�27/2021 A   ����DCSS_I�OC_T   �P $OPER�ATION  $L_TYPB7IDXBR1H[ �S2]2Rs�$�$CLASS  �������Pz��P� VERS?��  �1b�$' 2 ��P @ ���&8 J\n����� ���/"/4/F/X/ j/|/�/�/�/�/�/�/ �/??0?B?T?f?x? �?�?�?�?�?�?�?O O,O>OPObOtO�O�O �O�O�O�O�O__(_ :_L_^_p_�_�_�_�_ �_�_�_ oo$o6oHo Zolo~o�o�o�o�o�o �o�o 2DVh�z�������_�C_CCL ?���  	A�ll param~��
Base��Pos./S�peed che�ck(�Safe �I/O connect�}R���� �2�D�V�SIi�@{�� � ��� �I� D�V�h���������ٟ ԟ���!��.�@�i� d�v���������Я�� ����A�<�N�`��� ������ѿ̿޿�� �&�8�a�\�nπϩ� �϶����������9� 4�F�X߁�|ߎߠ��� ���������0�Y� T�f�x��������݇O�����%�N�I� [�m������������� ����&!3Eni {������� FASe�� ������// +/=/f/a/s/�/�/�/ �/�/�/�/??>?9? K?]?�?�?�?�?�?�? �?�?OO#O5O^OYO kO}O�O�O�O�O�O�O�}N�  ��OD_ m_h_z_�_�_�_�_�_ �_�_
ooEo@oRodo �o�o�o�o�o�o�o�o *<e`r� �������_ �SIh���b��� ������ӏΏ���� �(�:�c�^�p����� ����ʟ�� ��;� 6�H�Z���~�����˯ Ưد��� �2�[� V�h�z�������¿� ���
�3�.�@�R�{� vψϚ��Ͼ������ ��*�S�N�`�rߛ� �ߨߺ��������+��&�1�P%_�W�SOFDI10�y�2�y�3��y�4��y�5$��y�6��y�7��y�8�G�3�E�W�n�{� �������������� /FSew�� �����+ =Ofs���� ���//'/>/K/ ]/o/�/�/�/�/�/�/ �/�/?#?5?G?^?k? }?�?�?�?�?�?�?�? OO6OCOUOgO~O�O �O�O�O�O�O�O__ -_?_V_c_u_�_�_�_ �_�_�_�_oo.o;o Mo_ovo�o�o�o�o�o �o�o%7N[ m������ ��&�3�E�W�n�{� ������ÏՏ���� �/�F�S�e�w����� ����֟�����+�H=�H�Z�Od�v�O~� ������� ������&�A�Q� c���������ԿϿ� ���)�;�d�_�q� �ϬϧϹ�������� �<�7�I�[߄�ߑ� ������������!� 3�\�W�i�{���� ���������4�/�A� S�|�w����������� ��+TOa s������� ,'9Kto� �����/�/ #/L/G/Y/k/�/�/�/ �/�/�/�/�/$??1? C?l?g?y?�?�?�?�? �?�?�?	OODO?OQO cO�O�O�O�O�O�O�O �O__)_;_d___q_ �_�_�_�_�_�_�_o�o<o7oIo[o�ox�S�I����VOFF~noFENCE�o?EXEMG�o�o��cNTED�OP�oqAUTOT��[s����aMCC|pC�SBP�
PO�SSPD_ENB��jCONF_O�K�~F_IPARG_CR�z�g����~��o�q_�o;��o��`'�DIS�|'C_�r_`��y 