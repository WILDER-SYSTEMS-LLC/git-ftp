��   6�A��*SYST�EM*��V9.3�0146 5/�27/2021 A   ����PM_CFG�_T   � �$NU( HNL�  $IOD�_KEEP?ER�R_SEV?DE_V_FLG?CG	�CT
SCAN_M�ULT?CH1_wENB>CH2��FW: ECK?B�IND_ADDR>�PARE3�e~�    ���i�2��  �&STAT- ?\ $BD(?�UPDATE_F�W?PMTK_D�BGLV>PMU�IUEXPI_V�ERS? $CU�Rt �$$CL�ASS  �S�����b��b��xION�  1�'/ �b � �!�//(/:/L/^/����/�/�/ �/�/�/�??*?<? N?`?k/�?�?�?�?�?0�?���:���A