��   !��A��*SYST�EM*��V9.3�0146 5/�27/2021 A   ����BIN_CF�G_T   X� 	$ENTRI�ES  $QW0FP?NG1FU1O2F2OPz �?CNETG  ��DHCP_CT�RL.  0 �7 ABLE? �$IPUS�RE�TRAT�$S�ETHOST� �?�DNSS*� 8�D�FAC�E_NUM? $�DBG_LEVE�L�OM_NAM�� !�<�*� D $PR�IMAR_IG �!$ALTERN�1�<WAIT_�TIA �� FTޒ @� LOsG_8	�CMO>�$DNLD_F�I:�SUBDI�RCAP�� q��8 . 4� �H�ADDRT�YP�H NGT1H�� �z +�LS�&$R�OBOT2PEEyR2� MASK4�MRU~OMGD�EV�r���P�INFO� �$$$X �R�CMT A�$| ��QSIZ�X�� TATU�SWMAILSE�RV $PLA�N� <$LIN><$CLU����<$TO�P$C�C�&FR�&�JE�C�!�%ENB �� ALAR�!BF�TP�/3�V8 }S��$VAR79�M ON,6��,6A7PPL,6PA� -5�B +7POR��#_|12ALERT�&��2URL }>�3ATTAC��0�ERR_THRO��3US�9�!�8R0CqH- YDMAXN�S_�1�1AMOD�2AI� o 2A�� (1APWD � � LA �0�N�D)ATRYsFDE�LA�C2@�'`AERcSI�1A�'RO�ICLK�HMt0�'� �XML+ \3SGF�RM�3T� XOU̩3Z G_��COP c1V�3Q�'C�2-5R_AU�� � XR�N1oUPDXPC�OU�!SFO ?2 
$V~Wo��@YACC�H�QS�NAE$UMMY1��W2??�RDM�*	� $DISܤjSMB�
 7T �	BCl@DC1I2AI&P6�EXPS�!�PA�R� `RANe@ g ��QCL�/ <(C�0��SPTM
U� PWaR�-hCfV!SMo l5��!�"!%�7Y�P�% 0��fR�0�eP� _DcLV�Dey SNoB3 
j�hX_!`~�#Z_INDE,C�_pOFF� ~URnyD��)t�   t �!NpMON��sD�.�rHOU�#EyA�v��q�v�q�vLOCAܗ Y$N�0H_[HE��PI"�/  d	`ARPh�&�1F�W_~ d�I!Fap;FA�D8�01#�HO_� �R�2P$`�S�TEL�	% P K � !�0WO�` �QE� LV�k�2H#ICE�ڀ����$d�  �S������
��
���`S$Q��  1b�$'�0 �
���F��p��"�S�L��$� 24�����@��e��� 4���! �0ʟ����-�4�Ɵ ��8�I�L���p_V`4��S�z��� ����¯ԯ���
���.�@��� _FLT�R  �?� *��������ޛndx4�2ޛ8�SHE`�D 14� P'��I�ٿ��:� ��^�!ς�Eώ�iϷ� �ϟ� ���$���H�� l�/�Aߢ�e��߉��� �������D��h�+� ��O��s������
� ��.���R��^�9��� ��o����������� <��r5�Y� }����8� \�Cy�������PPP_L��A1e�x!1E.9"0/�8%1I/>�255.�%@/&��Q�7#2>/P.@� d/v/�/�/�&3�/�P.-0�/�/ ??�&4 .?P.�0T?f?x?�?�&5�?P.@�?�?�?O�&6OP.�@DOVOhO�zOT�aP��0���8(�Ӱ��� Q�	 ��N<0_e_w_J_��_�_�_�_�_�_�P �_%o7oIoomoo�o@�obo�o�o�o�N�o�T�5 |
ZD�T Status��oD����}�iRConnec�t: irc�t/?/alertb~� ��+��wtY�k�}�P�������A�d�RJ������ ��$� 6�H�Z�l�~��������ƟQs$$c962�b37a-1ac�0-eb2a-f�1c7-8c6e�b555bb26  (H��l=�O�Ha�s���A��X�'R��)z��P��*s,P!T,$4�񯨰*! ߯��@�'�M�v�]� ������п����ۿπ���N�5�r�Y��棧�&%PDM_�Q	&+"SMB 
&%U�#l��O����� I߿�ś�����_CLNT 2&)9�4+t	�|�#| j߯ߎߠ�������� ���Q�0�u��f�������
.SMTP�_CTRL R� P%��4�	t��"� c���R���v���#|��	N�Q�΢��=7����� S���USTOM ����&P |�TTCPIP���'xU"Ri E�L$&%#Q� H�!TP	��?rj3_tpт���+ ��!KCL��������!C�RT.uR�?!CONSv�
��ib_smo	n~r