��   (�A��*SYST�EM*��V9.3�0146 5/�27/2021 A 	  ����PASSNA�ME_T   �0 $+ �$'WORD � ? LEVEL � $TI- OUTT�&F/�� $SE�TUPJPROG�RAMJINST�ALLJY  $CURR_OަUSER�NU�M�STSTOP�_TPCHG �V LOG_P NT��N�  6 C�OUNT_DOW�N�$ENB_�PCMPWD� �$DV_� IN�� $C� CR5E��A RM9� =T9DIAG9(|�LVCHK >FULLM/��YXT�CNTD��MENU�A�UTO+�FG_wDSP�RLS��U�BURYBA�N��GI�  �&ENC/ � CRYPT�E ���$�$CL(   ���[!�� d P �V� IONX(�K 1b�$D�CS_COD?����_%�  W�'_� �/�(S  JZ*�� \ �&�A�91�"[!	? 
 $b!�� =?4?B?X?f?|?�? �?�?�?�?�?�?OO�0O>OTOL#'SUP
�  :�VOhO�#F��O�O�O�� � \Q��_ �0�� V�[_t&��j���D�Op_��.W,_��K!��U�_oKLUGH �1[) K �)�_oo/oAo Soeowo�o�o�o�o�o �'�_�o#5GY k}������o ���1�C�U�g�y� ��������ӏ��	� �-�?�Q�c�u����� ����ϟ�����)� ;�M�_�q��������� ˯ݯ���%�7�I� [�m��������ǿٿ ����!�3�E�W�i� {ύϟϱ��������� ��/�A�S�e�w߉� �߭߿��������� +�=�O�a�s���� �������� ��'�9� K�]�o����������� �������#5GY k}������ ��%