��   !�A��*SYST�EM*��V9.3�0146 5/�27/2021 A   ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_  �$$�CLASS  O�����D���DVERSIO�N  �1b�8LOO�R G��DD<Z$?���q���M,  1 <DYX< [�����D'�i���B��i!/W/ �@��C/e/�/y/_ �"�/�/�(�$M�NU>A>"��� n <�&�U�����7���"?��;1I��;��|�1J��E0D�X�^���a�����=7���%����-<&+��?�z;S�;�s���m�E0�D�'������o�u9;��^}���:�E��E0u;�H�v�a>;`�߶:KG�U0����)[�-D��לo��%���<�>�?��ؼ�T��0��<9�g�<Lg�<<�?�Q��L�'�R��� �%�8��<��A�@(=���Wſ�<�8���<}<�<��@P�M����=Ӆ�!R�)O;EV�E@&<�8#h�<�k<�;��@Z�8�)}H�!N�)�5@�9@ܼ@�G�A@i�Dc�="j�<;�@S�N���G��!��J�)��W%��~�>;�u*?�~|���<�������;��@�RD����6ȇ�_�!��9E?W?i4\q?'_ 9_k?]_o_�_�_�_�_ �_�_�_�_o#o5ow7�<d�����<���?ۄ�<lCX<�g���QD<��@��:D��tC7?A��`z.�<8ʃ2�4��?�0�����F��`�EoWoio{o)�;M_u<��%��<���<&	���`{;�
;�#f�3�}p��D	�0L�>?�~�D<Ϥ=���a�*�?��x<�\����}�ч�?�~�GD+�(�cO�đ��u9�=�C�}J����8?|��=�Eڻt;��;x_>�f����p�Ċ*��9�۲Ï�����uw��o�Z=�:�r�@�g�����?<�{	?���D!��a����eju;���;zȃ=|����?�?����p1W�|�B�<lƃ=�/D$����a�V�j�$�u:{�w����C�4��:���H�p�;�:�>4�ݻ'JQ��[D!K;�a����DZ�u:h���<�@>տ=Q�e�qm�l������p#�=%\?h��D>�+�b��Ęw�u;��;����=j�����?�μ�LS��jUU<�F��?��D�%)��bOL��mdAx6�z�7�>LS=Fdy�>K�?zݤ��8��K�*���g4����D���e���T9�u:Q���<��3����<*�L?���=5��?����-K�?Q||�D2"�aE��*~�u:|g�;+��>4+#�:Ξ	P}���D��4.g<���-?{��D&����b">�y�"�ً�����оG��;����p(;���>G�x��0M����_�a����A�Ku;�G����<�7m;����0u�4E����P<5eg�?��D"Q��a�\�c�	�u;�ؼ.A=Փ<!/}@�ļK���V��<Q�:?���D��ae�%�h�u:z[���K+G�Um�<B��������>Uv':���_?z`1D���a1��$�Zu:f>���)�����<�&���`\�4���>�����r?fB2D3����a�ák�'����:di����u�b���y���;����:�ލp��Č���=��Ï��a��/�� ����Ͽ����3���K�i�O��6|����4=�G(��l�?}�q��r~��a���s���E��x��P4�c/u:z��ώ������ ��Y��6��??�3���
ڍ��=�>���Խ#|��?X�D�����aI��V ��3ߝ�Gߥ��߹����v�e;8��>��6�;�
�?�����
���0=`m?�v�D(��bR�Ă
�u:�1��=oV?�87K<���?�l��sϿ�8U�=p��?�1D`�v�?d�Uħ;�q����ߐ���o�ݺ�H}��ǿ;;����2�-%>���@��%c?o��D+wT�a�vF���Ax8��]:�#�= �ߒ����0,��F0�� �<�E^�?ȤD�$��ao���i/��{����f>2݊;5�n)@м��2��<����?|kD)$��a��ĉ����{���"Խ�9�:��V�0�)�F,=�E��<B��?~���D!p�a��c�7�@�{��;1��=�m���w��`T�*�����y�<'��F?~��D'�;���n�~Þ y��������+# EsY{���� ���'/]C e�y����� /�/G/-/?/a/�/ u/�/�/�/�/�/�/�/ ?C?)?K?y?_?�?�? �?�?�?�?�?�?-OO 5OcOIO[O}O�O�O�O �O�O�O_�O_1___�EZ�z��|���:�R;�7��m�.�U�W=:���<P�S?��fD����?�>�P����g_ �_{_�_o�_�_!oOo 5oWo�oko�o�o�o�o �o�o9Ao Ug������ �#�	��=�k�Q�s� ������׏��Ϗ�� �'�U�;�]���q��� ��ӟ��۟	���?� %�7�Y���m��������ů�ٯ��;��[��~;A*��*?߉�@�	���:��;*����������D0��]�cɴ�Y���_C���W����ɿ ۿ��+��3�a�G�i����}Ϗϱ������$�MNUFRAME�NUM  ������D � �4�T�OOL A����6��� � <����_���'	?��3;�.c�c�����dѓ՟�o��z?��C���ɟհ�ٓѓՏ�B��Ж?ٚA�33�������A��Љ��A������A��Й�L�B��8�J�����dз�q����?�B��������d������� ���7� ��/���c߭�wߥ��� ������+3aG@Y{��/���
	
 