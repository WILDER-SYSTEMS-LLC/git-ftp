��  Ij�A��*SYST�EM*��V9.3�0146 5/�27/2021 A   ����SBR_T �  | 	$S�VMTR_ID � $ROBO�T9$GRP�_NUM<AXIaSQ6K 6NFF�3 _PARAM�F	$�  �,$MD SPD�_LIT  &2j*� � �����$$CLASS  ���������� VER�SION��  1b�$�'  1 � �T���R-�2000iC/2�10L���  �aiSR30/}3' 160A���
H1 DSP�1-S1��	P�02.009, � 	�  �  ��  �!��  8�w���������
=��9�9~��	d���� ��� ,��� � sW�� ����< RR���  ������  2>,���>�����
��ߠ	/���&������o�� T���w�����_� �<���`�?���~ ���:c	`�D 0 ���� g� :�?��:~}'bx�E/�/�/�/�/����/��3?C?U?�Z�r?�?�?�?�?����0�D40/4LY2�^2fx����������������a��w���9 :�� @m�B�|��݊���8��8������� 4�����<]�i�A�_	�+��,  +��4 C8$y�?R$���\'��
�����!�G5"B	�� � 2 �tB� ��#9=�"��	-�Ou_0�_�_�_3а_ ? �_�_oo1oCoUogoyo�?�? �2HO�H3^�R"O4O�����PA��~VO��nJ�8H~@�C0r�$� o ��/G�G��M����2�%_
 &����:s0��y�+� � ���� ��T��zo���ƻ�3X��:�r���"*W �6SU�>PS"S �	�zLTOTY���`-�?�Q�c�3	�h� �_����ŏ׏������1��o�o �2RU1�d4	I4^4�o��m�=���(���sq�rp@ ?~��%/nB2�� 0���  ���ύ��"Ls$@���}#�5����@��pK8$�E�������\'
��}U����؍���~! f s< ��q�u�#����
,��� >q������4
( ���f F�k�}�������ſ׿��D�V� j�T5b^5�������pƟ�؟������q�!����� W��pJ8$��Ͼ���\ )�����F�+�՚�� ����ʯܯ�߷���$� ��H���#�5�G�Y�k�`}������ "�
T6^6F�X�j�TO�Ϣ�����s���ϟ������)�p�4 � :"o|��x"���\'���i	��0/
�ꚨ�^�p� �ߔ�]o��ߐ � ����#5G�Y��>�EX�TENDED AsXI���7�0�8�c8	F��H rA cT�0.3����� P��FB&�����z ��ߟ�  {��H�?�Su%��03sARR��
O �0/ B/T/f/x/�/�/�/����t� d �A �c A��:TY:q�/?? 1?C?��a?s?�?�?��?�?�?�?�?O�\�?����OH('@&O��KL	KH�E@�O�O�O�O�O�O �O__&_8_J_\_n_��_�_�_�_�_�_�\� �_o o2oDoVohozo �o�o�o�o�cDO6O�o ZOlO~OFXj|� �������� 0�B�T�f�x������_ ��ҏ�����,�>� P�b�t��o�o�� *���(�:�L�^� p���������ʯܯ�  ��$�6�H���Z�~� ������ƿؿ����  �2ώ�W�J�ğ֟� ����������
��.� @�R�d�v߈ߚ߬߾� �������b�*�<�N� `�r��������� ��l�^���ϔϦ�n� ���������������� "4FXj|� ��� ��� 0BTfx���� *���@�R�/,/>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?��?�?�?�?�?�?  OO$O6OHOZO�O rO��/�O�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o �?Rodovo�o�o�o�o �o�o�o�O�O0 �O�O�O����� ���&�8�J�\�n� ��������ȏڏ�Ho �"�4�F�X�j�|��� ����ğ RD�h zB�T�f�x������� ��ү�����,�>� P�b�t�����􏪿ο ����(�:�L�^� pς�ޟ�Ϛ��&�8�  ��$�6�H�Z�l�~� �ߢߴ����������  �2�D�Vﲿz��� ����������
��.� @��Ϯ�X������Ͼ� ������*<N `r������ �p�8J\n �������H� z�l�5/����j/|/�/ �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?OO,O>O PObOtO�O�O�O/�O �O</N/`/(_:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o �?�o�o�o�o�o�o  2DVh�O�O� �O__��
��.� @�R�d�v��������� Џ����*�<��o `�r���������̟ޟ ���p��]�� �������ȯگ��� �"�4�F�X�j�|��� ����Ŀֿ�D���� 0�B�T�f�xϊϜϮ� ����.�����d�v��� P�b�t߆ߘߪ߼��� ������(�:�L�^� p�����������  ��$�6�H�Z�l�~� ����Ϩ�"�4�F�  2DVhz�� �����
. @Rd����� ���//*/</�� �����/�����/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? Ol"OFOXOjO|O�O �O�O�O�O�O�OV/_ _�/�/�/x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o *O�o(:L^ p����4_&_� J_\_n_6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z����o ��ԟ���
��.� @�R�d������� ������*�<�N� `�r���������̿޿ ���&�8ϔ�J�n� �ϒϤ϶��������� �"�~�G�:ߴ�Ưد �߲����������� 0�B�T�f�x���� ��������R��,�>� P�b�t����������� ��\�N���r߄ߖ�^ p�������  $6HZl~ �������/  /2/D/V/h/z/�/�� �/0B
??.? @?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `O�rO�O�O�O�O�O �O__&_8_J_�/o_ b_�/�/ ?�_�_�_�_ o"o4oFoXojo|o�o �o�o�o�o�o�o zOBTfx��� ������_v_ � �_�_�_��������Ώ �����(�:�L�^� p���������ʟܟ8  ��$�6�H�Z�l�~� �������B�4���X� j�2�D�V�h�z����� ��¿Կ���
��.� @�R�d�vψ�䟚Ͼ� ��������*�<�N� `�r�ί�ߊ���(� ����&�8�J�\�n� ������������� �"�4�F���j�|��� ������������ 0�ߞ�H�����߮ ����,> Pbt����� ��/`�(/:/L/^/ p/�/�/�/�/�/�/8 j\%?��Z?l?~? �?�?�?�?�?�?�?O  O2ODOVOhOzO�O�O �O/�O�O�O
__._ @_R_d_v_�_�_�/�_ �_,?>?P?o*o<oNo `oro�o�o�o�o�o�o �o&8J\n �O������� �"�4�F�X��_�_p� �_�_o֏����� 0�B�T�f�x������� ��ҟ�����,�� P�b�t���������ί ���`�����M��� ����������ʿܿ�  ��$�6�H�Z�l�~� �Ϣϴ�����4����  �2�D�V�h�zߌߞ� ���������T�f�x� @�R�d�v����� ��������*�<�N� `�r������Ϻ����� ��&8J\n ����ߘ�$�6�� "4FXj|� ������// 0/B/T/��x/�/�/�/ �/�/�/�/??,?� ��u?���?�?�? �?�?OO(O:OLO^O pO�O�O�O�O�O�O�O  _\/_6_H_Z_l_~_ �_�_�_�_�_�_F?o o|?�?�?hozo�o�o �o�o�o�o�o
. @Rdv���� _����*�<�N� `�r�������$oo�� :oLo^o&�8�J�\�n� ��������ȟڟ��� �"�4�F�X�j�|�� ����į֯����� 0�B�T����ԏ���� 
�ҿ�����,�>� P�b�tφϘϪϼ��� ������(߄�:�^� p߂ߔߦ߸�������  ��n�7�*錄��ȿ �������������  �2�D�V�h�z����� ��������B�
. @Rdv���� �L�>��b�t��N `r������ �//&/8/J/\/n/ �/�/�/ �/�/�/�/ ?"?4?F?X?j?|?� 
��? 2�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_�/b_�_�_�_�_�_ �_�_oo(o:o�?_o Ro�?�?�?�o�o�o�o  $6HZl~ �������� j_2�D�V�h�z����� ��ԏ���tofo� �o�o�ov��������� П�����*�<�N� `�r���������̯(� ���&�8�J�\�n� ������ �2�$��H� Z�"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�x�ԯ�߮� ����������,�>� P�b﾿��z����� ������(�:�L�^� p���������������  $6��Zl~ �������  ���8������ �����
//./ @/R/d/v/�/�/�/�/ �/�/�/P?*?<?N? `?r?�?�?�?�?�?( ZLOp�JO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�/�_�_�_�_oo 0oBoTofoxo�o�?�o �oO.O@O,> Pbt����� ����(�:�L�^� �_��������ʏ܏�  ��$�6�H��o�o`� �o�o�oƟ؟����  �2�D�V�h�z����� ��¯ԯ���
��x� @�R�d�v��������� п���P���t�=Ϙ� ��rτϖϨϺ����� ����&�8�J�\�n� �ߒߤ߶���$����� �"�4�F�X�j�|�� ��������D�V�h� 0�B�T�f�x������� ��������,> Pbt��ߪ�� ��(:L^ p������&��  //$/6/H/Z/l/~/ �/�/�/�/�/�/�/?  ?2?D?�h?z?�?�? �?�?�?�?�?
OOx ��eO���O�O�O �O�O�O__*_<_N_ `_r_�_�_�_�_�_�_ �_L?o&o8oJo\ono �o�o�o�o�o�o6O�o �olO~O�OXj|� �������� 0�B�T�f�x������� 
oҏ�����,�>� P�b�t������� *<N�(�:�L�^� p���������ʯܯ�  ��$�6�H�Z�l�ȏ ������ƿؿ����  �2�DϠ�ҟğ��� ����������
��.� @�R�d�v߈ߚ߬߾� ��������t�*�N� `�r��������� ���^�'���Ϧϸ� ���������������� "4FXj|� ����2�� 0BTfx��� �<�.��R�d�v�>/ P/b/t/�/�/�/�/�/ �/�/??(?:?L?^? p?�?�?��?�?�?�?  OO$O6OHOZOlO� ���O/"/�O�O_  _2_D_V_h_z_�_�_ �_�_�_�_�_
oo.o @o�?Rovo�o�o�o�o �o�o�o*�OO B�O�O�O���� ���&�8�J�\�n� ��������ȏڏ��� Zo"�4�F�X�j�|��� ����ğ֟�dV � z��f�x������� ��ү�����,�>� P�b�t���������� ����(�:�L�^� pςϔ��"����8� J��$�6�H�Z�l�~� �ߢߴ����������  �2�D�V�h�Ŀz�� ����������
��.� @�R���w�j������ ������*<N `r������ �&��J\n �������� /��~�(/�������/ �/�/�/�/�/�/?? 0?B?T?f?x?�?�?�? �?�?�?@OO,O>O PObOtO�O�O�O�O/ J/</_`/r/:_L_^_ p_�_�_�_�_�_�_�_  oo$o6oHoZolo~o �o�?�o�o�o�o�o  2DVhz�O� �__0_�
��.� @�R�d�v��������� Џ����*�<�N� �or���������̟ޟ ���&�8���P� �����ȯگ��� �"�4�F�X�j�|��� ����Ŀֿ����h� 0�B�T�f�xϊϜϮ� ������@�r�d�-߈� ��b�t߆ߘߪ߼��� ������(�:�L�^� p����������  ��$�6�H�Z�l�~� ����������4�F�X�  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/����x/���/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4O�XOjO|O�O �O�O�O�O�O�O_h/ �/�/U_�/�/�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o<O�o(:L^ p�����&_� �\_n_�_H�Z�l�~� ������Ə؏����  �2�D�V�h�z����� �oԟ���
��.� @�R�d�v������� �,�>���*�<�N� `�r���������̿޿ ���&�8�J�\ϸ� �ϒϤ϶��������� �"�4ߐ�¯��}�د ꯲����������� 0�B�T�f�x���� ���������d��>� P�b�t����������� ����N�
�ߖߨ� p�������  $6HZl~ ����"���/  /2/D/V/h/z/�/�/ �/,�/BTf.? @?R?d?v?�?�?�?�? �?�?�?OO*O<ONO `OrO�O��O�O�O�O �O__&_8_J_\_�+��$SBR2 1��%�P T0 � ���/�' �_�_�_�_oo &o8oJo\ono�o�o�o�o�Q��o�_�o '9K]o��� ����o��o#�5� G�Y�k�}�������ŏ ׏�����z��� Q�c�u���������ϟ ����)�;��_� B���������˯ݯ� ��%�7�I�[�m�P� ��t���ǿٿ���� !�3�E�W�i�{ύϟ��x�Ϡ������� )�;�M�_�q߃ߕߧ������{~i_���!� 3�E�W�i�{���� �����������(�:� L�^�p����������� ���� $��Z l~������ � 2DV:L �������
/ /./@/R/d/v/�/l �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �/�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�?_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo_BoTofoxo�o �o�o�o�o�o�o ,>P4ot��� ������(�:� L�^�p���f����ʏ ܏� ��$�6�H�Z� l�~���������؟� ��� �2�D�V�h�z� ������¯ԯ��ʟ
� �.�@�R�d�v����� ����п������� <�N�`�rτϖϨϺ� ��������&�8�� F�n߀ߒߤ߶����� �����"�4�F�X�j� Nߎ����������� ��0�B�T�f�x��� ������������ ,>Pbt��� �����(: L^p����� �� /�$/6/H/Z/ l/~/�/�/�/�/�/�/ �/? ?2?/V?h?z? �?�?�?�?�?�?�?
O O.O@OROdOH?�O�O �O�O�O�O�O__*_ <_N_`_r_�_hOzO�_ �_�_�_oo&o8oJo \ono�o�o�o�o�_�_ �o�o"4FXj |�������o ��0�B�T�f�x��� ������ҏ����� �>�P�b�t������� ��Ο�����(�:� L�0�p���������ʯ ܯ� ��$�6�H�Z� l�~�b�����ƿؿ� ��� �2�D�V�h�z� �Ϟϰϔ�������
� �.�@�R�d�v߈ߚ� �߾���������*� <�N�`�r����� ����������8�J� \�n������������� ����"4�*�j |������� 0BTfJ\ ������// ,/>/P/b/t/�/�/| �/�/�/�/??(?:? L?^?p?�?�?�?�?�? �/�? OO$O6OHOZO lO~O�O�O�O�O�O�O �O�? _2_D_V_h_z_ �_�_�_�_�_�_�_
o o.o_Rodovo�o�o �o�o�o�o�o* <N`Do���� �����&�8�J� \�n�����v��ȏڏ ����"�4�F�X�j� |�������ğ����� ��0�B�T�f�x��� ������ү�ȟڟ� ,�>�P�b�t������� ��ο������� L�^�pςϔϦϸ��� ���� ��$�6�H�,� V�~ߐߢߴ������� ��� �2�D�V�h�z� ^ߞ����������
� �.�@�R�d�v����� ����������* <N`r���� ����&8J \n������ ��/�4/F/X/j/ |/�/�/�/�/�/�/�/ ??0?B?&/f?x?�? �?�?�?�?�?�?OO ,O>OPObOtOX?�O�O �O�O�O�O__(_:_ L_^_p_�_�_xO�O�_ �_�_ oo$o6oHoZo lo~o�o�o�o�o�_�_ �o 2DVhz ��������o �.�@�R�d�v����� ����Џ����*� �N�`�r��������� ̟ޟ���&�8�J� \�@���������ȯگ ����"�4�F�X�j� |���r���Ŀֿ��� ��0�B�T�f�xϊ� �Ϯ��Ϥ������� ,�>�P�b�t߆ߘߪ� �����������(�:� L�^�p������� ���� ��$��H�Z� l�~������������� �� 2D(�:�z �������
 .@RdvZl �����//*/ </N/`/r/�/�/�/� �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �/�?O"O4OFOXOjO |O�O�O�O�O�O�O�O _�?0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>o"_boto�o�o�o �o�o�o�o(: L^pTo���� �� ��$�6�H�Z� l�~������Ə؏� ��� �2�D�V�h�z� ������ԟ����
� �.�@�R�d�v����� ����Я���؟�*� <�N�`�r��������� ̿޿���&�
�� \�nπϒϤ϶����� �����"�4�F�X�<� fߎߠ߲��������� ��0�B�T�f�x�� n߮����������� ,�>�P�b�t������� ��������(: L^p����� ����$6HZ l~������ �/ /D/V/h/z/ �/�/�/�/�/�/�/
? ?.?@?R?6/v?�?�? �?�?�?�?�?OO*O <ONO`OrO�Oh?�O�O �O�O�O__&_8_J_ \_n_�_�_�_�O�O�_ �_�_o"o4oFoXojo |o�o�o�o�o�o�_�_ 0BTfx� ��������o �>�P�b�t������� ��Ώ�����(�:� L�