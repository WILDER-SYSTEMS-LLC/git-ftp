��   ��A��*SYST�EM*��V9.3�0146 5/�27/2021 A 	  ����DRYRUN�_T  4 �$'ENB � $NUM_P�ORTA ESU�@$STATE� P TCOL_���PMPMCmGRP_MASKZ}E� OTIONN�LOG_INFO�NiAVcFLTR_EMPTYd $PROD__ �L �ESTOP_�DSBLAPOW�_RECOVAO{PR�SAW_� �G %$IN�IT	RESUM�E_TYPEND�IST_DIFF>A $ORN41p� d =RVR &�J_  4 �$(F3IDX؞�_ICI ��MIX_BG�-y
_NAM�c MODc_U�Sd�IFY_T�I� ��MK�R-  $�LINc   �"_SIZc?��� �. h �$USE_FL�C 3!�:&iF*S�IMA7#QC#QB�n'SCAN�AX֋+IN�*I��_C7OUNrRO( ���!_TMR_VA�g#h>� ia �'` �����1�+WAR�$ҵH�!�#N3CH��PE�$O�!PER�'Ioq7iOq� ���OoAT�H- P $ENABL+��0BT���$$CLASS ? ���A���5��5�0VERS��G  �1b�6/ E�5�������-@]F@AbE���%A�O���O�O��X��3EI2>K�0 __0_B_T_f_x_�_ �_�_�_�_�_�_oo0,o�O*W?"HI@ ��lo��V0.|j�|m�� �� 2>I  �4%DATAM�AP:o�� qT��%OFFSEOSI�� �o��h�$J%PL�C!ET%( �RU>�%Y�	bAqoAt�� ���f����R�1���c$"+ �ktK-@�����bA��X lA-@vNڏ��� �"�4�F�X�j�|��� �����{[EoAǁoA� ��
��.�@�R�d�v����������ЯDZLax R�cC!2�lǏ1�C�U�g�y� ��������ӿ���	� Ɯ#�<�N�`�rτϖ� �Ϻ���������� 8�J�\�n߀ߒߤ߶� ���������"�-�F� X�j�|�������� ������)�;�T�f� x��������������� ,7�Pbt� ������ (:E^p��� ���� //$/6/ ASl/~/�/�/�/�/ �/�/�/? ?2?D?Ch �4�0��{?@