��   #��A��*SYST�EM*��V9.3�0146 5/�27/2021 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	  /GR�P: $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2(��� RING��<�$]_d�REL�3� 1 N ��CLo: �� �AX{  o$PS_�TI����TIME z�J� _CMD���"FB�VS �&C�L_OV�� FR�MZ�$DEDXv�$NA� %�OCURL�W����TCK5�F�MSV�M_LIF	��;8�G:w$�A9_0M:_ ��=�93x6W� �">�PCCOM���FB� M�0�MAL_�ECI��PL!�"DTYkR�_�"�5L#�1END�D��o1 e�5M�P PL� �W �  $S�TAL#TRQ_MH��0KN}FS� ��HY�J� |GI�JI2�JI�E#3AnCuB��A� �$�AS=S> ���	Q������@VERS�I� W � 1b�$S �1'X ���N ��n_Y_��_}U����q��� ����%�	?��Lu_�_��_�Q�pߎ�����
�� B�!�1<�\2P+f���,m�UQToT�V$���������g�c�N��K��F����_�o�\lg�o�o�o��ox� 7q�z=p$�eB@Mu @
BZpYqYq@�_z#w���d�p�����=L̔g�%���?�/���@� O�t���������Ώ������(�:�� �	Ue�s�]���T  2�ğ֟����� 0�B�T�f�8b���� ����Ưد���� � 2�D�V�h�z������� ¿Կ���
��.�@� R�d�vψϚϬϾ��� ������*�<�N�`� r߄ߖߨߺ������� ��&�8�J�\�n�������<������� ��&�8�J�\�n������|(�������� ��2/hS��w�����
��$&4 1D\���O���K1���L�.O���O!�6Q�A���H��L��	�L5uD��;Eq��B�{@\�C�� ��B�� ���B6�?��XRUB����B�B)B9�Mǡ���	I�P�^M�>�L��wF�X�G?��C��b�� �A�  /�>��F2J[�U�*���g/��/v/�/�+��T�'U5#Y&�$N@ ^��&�Q� � ��U/�6"�?��B���¶��˹Bm�B��G��%�����B��#��`x��I�B��B����FB��)>�)��?�,�@*(�־\��?z�>o�WB��� �]�%JO�B_DBL_SA�D@68�/Y�� "�\�1��!�5���B4��h���B�0�δ�t!_ġ�O��)�0�B4����0�0s��8�t"�=9��� �DD@��->z :�����:���׾B�  Ԏ2�not a program�?�TQ��4F��!��_��B�?��$2��B�65Bs6��B)Ĵ�p��)��X�B�9_�$�@�@���@p�M<;� �>ޕ�@C�:���	�>��6��)8N2P'�2�ROS_MOVE�SM_WILDE�RnO[�X��1P���2�B����B�/�"B��B�R���@i�:��B��^eB��-�B��bBיKNj]��@�%���@���I��4>��X>	#�!b�I@__�0_BX�vS�{B����%B��,wB��[B�kH��@hn[�`���HB�+_�B��W&`�@�e�);���5��@��h�X�پ>ٶ��T�s�:O�_�_�_BX��vS��B�����
^B�.IB���B�\��@�dn[�B���`�BĿ�RB�S��@c��Z�d`(��@��A�KX>�'+>1�b��o�o��o?[�vS�B��<��F`r�B���B�N��}�pFB�������F`8B��_�B�Q �@`�)�:�Q6�@�R��[�r>�U��@�{;I[m�Y�1�m�!@���RB�x���B��7����&b�@@��)@�^�B�p����B�_�	�9��'W�`j���x�?x�&�@>���A��@��@��N.�;K��S�CI_TAI�0W�ITCH+�xE GaKB�T#�a�U������U�@0���������B9�Ъ@1�)�#A��@�]P����>��&�7@�{;
�fҏ��yD�]wF�Sf���!�"!@��t��@�eBK�MfBrS�Bl?N�ċL͞)Ґ�)@�3�@��aBKY�BrD_Bl/Vꐁ�)��ާ����!�@�ɿ��?fB�?${��<<��|m�%CLAMP��j�I@{��BUTK�HvR�@vAޔ	���
B��PB���B�=���Н*�@8lA���¨��B��w�B�Bׯ�ͪ��)���@1P�>;��*?q�@�?��?��=qL�`��?�082k�xE� ���S� Y;vR���A��&�n�L��gB���DB�tġ��jnZ�-A��{	�nV
��B��bB�Cġ���)?�I���~_�@���?�l�=���ȿm�7%x���� ��2���TZ͒�)��Ak$|¦���B2qxB���(B�GQĶ� �)�AAj�_¦v��"��s&��*�/Vn-��@�˪�+��#>��Z��T������L��ϾsJ ���5T�a3�v��}A����n.#��YB���B��t�0�n���A�(�m�K���qB��,B��O�� =+b�����@@�x+�>��g>��ȟ���w:;K�`��βUF_RI�VETLOCAT'ION��yD W� ��=�N��R�@�����%����_B��MB��h���n���lu@�;�����f��@�B���B������sn�4����$G@�<���?jQ�?�9�Bd�����P�b�t߆ԭN��{�>@�����foB��B?��9��A�s���ze@����W���^�!b�Bf��4j��z#qIx�@�<�=��p������#;{;���SO��pM����Kv��	 l>�n�{�3B��;B�MN�ϻ��A�-%�nP����B��B�N�*�;��� �z8@���;>�
�>�?ٰ��M���L��TOOL_2_�PICK_APR�OA��zC>YT���n�p��A���a �ABD�@�B�S�B��SĶ��p���A��� �o�BDBlB�?N�B�@����q����@t�y�����?�t��?Q�Gz<
  cX��_�z�����r���)A�{�� e&BDD�B�R\B�?��������|A��v� c@BD�C�B�W]� E�����-�B3@���нWZ�>𗙻7@qLI�m�B��&W�vR�_yA-�x��}[r6K�B�tzB���Ġ�qnZ��G�A-=��}g��w�B��>�B�rĠ�V������rR��@��w?�52��ߞ.�>4�A������ο_�57+���!���
/�CyD�$PL�CL_GRP 1�ǐ��;!��~ �A��|0T*m?p?h�ET)�/ �/�	�/�/�/�/�/? �/%??I?4?m??N,�n�T"h=?nAl)