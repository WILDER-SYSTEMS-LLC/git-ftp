��   v��A��*SYST�EM*��V9.3�0146 5/�27/2021 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@ � &�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	� �&USRVI| 1  < `��R*�R��QPRIƍm� t1�PTR�IP�"m�$$C�LASP ��)�a��R��R `\ �SI�	g  1b�$'�2 ���R	� ,��d?���aa1`jb�ed`a����? � �`dc<�o��
 ��a�o@�o�o%7 �o \n����E� ���"�4��X�j� |�������ďS���� ��0�B�яf�x��� ������O������ ,�>�P�ߟt������� ��ί]����(�:� L�ۯp���������ʿ�ܿa`TPT�X��l����a`� s縄�$/s�oftpart/�genlink?�help=/md�/tpmenu.dg޿xϊϜϮ�g� ��������,߻�P� b�t߆ߘߪ�9߻��� ����(�:���^�p�`��������a��f�b��g ($R������6�!�Z���4`ada��c������� N��k
$��aJ��aJ� � �J�	H���E���跪����b���`  ���H G�p��J#�J�Ffbc :c�B �1)hR �\��_�� wREG VED?����wholemod.htm�	�singl�d�oubtr�ipbrows3b�i{� W�����"/�����dev.s��lo/� 1r,	t�/A�//K/�/�/ ?�/5?G?Y?k?}?�?� ��?�?�?�? OO+O=OOOaOjE2P �?�O�OqO�O�O�O�E �	�?�?_/_A_S_e_ w_�_�_�_�_�_�_�_ oo+o=oOoao/'yo so�o�o�o�o�o�o 1CUgy�� �����? �2�D� V�h�z��������O ���Ǐُ.�@��O	_ ���������П˟ݟ ���%�7�`�[�m� ��������oկϯ�� �!�3�E�W�i�{��� ����ÿտ����� /�A��|ώϠϲ��� ���������B�T� #�5ߊߜ�S�e�K��� �����,�'�9�K�t� o���������� ���߯1�+�Y�k�}� �������������� 1CUgy�� k���� 2D Vhzuߞ�� �����ߧ@/;/M/ _/�/�/�/�/�/�/�/ �/??%?7?`?[?m? ;��?�?�?�?�?�?�? O!O3OEOWOiO{O�O �O�O�O�O�O�O�4_ F_X_j_|_�_�_�_�_ �_��_o�_�_BoTo�bj�$UI_TO�PMENU 1�-`�aR� 
d�aQ)�*default�_ ]*lev�el0 *[	 #�o�0�o�o�o�	rtpio[23�]�8tpst[1=xY�o�o�=�h58e01_�l.png��6menu5�y�p�qC13�z�r�z�t4�{��q��?�f�x��� ������RT�������1�C�҄pri�m=�qpage,?1422,1J��� ������˟֏����%�7�I�ؖ^�class,5R�����Ы���ϯڔf�13�֯��0�B�T�ۓ^�53p�������ƿؿۓ^�8��%� 7�I�[�ڟϑϣϵ�����Y�`�a�o߀�mΙq�;�mCvt�yN}6Hqmf[0�PN�	��c[164=w��59=x�q)�L[��tc8�|�r2� �}Q����w�{��O� ������ ��$�o� H�Z�l�~�����Q�c�80������	-`�r�22gy�� �>p���	- ����n����e�w�1���//*/�</7�^�ainedi	�s/�/�/�/�/�2�config�=single&>^�wintpj��/ ??*?<?����r?!�>��gl[57�ٕ Sߵ?�;Ip�08�ݔ0A7�9�?�6���62,O[6�:�?OqO�x�6�z�4s�x�O ���x� �B�Q�*_<_ N_`_r_�_3��_�_�_ �_�_o�_&o8oJo\o�no�o�o�!;�$dokub�%oc�13~��&dual�i38���,4�o�o�o9 �o�n�o�ax�� #o�������%�3.=_!g�Q�b8 "�z�������\ԏ提��
���+:6��i48,2Q��b]������ ]?ҟ�/�UE߻����s���_����G�u��:���"�f7.�ݣB�Or��J�\�6G�u7������ÿտ翮��27��)�;�M�_�q� � �U�����������!�1�/�A�S�e� wߪ�߭߿������� ���+�=�O�a�s�� ���������������6
�?�Q�c�u����$��74�����������C���6�	�TPTX[209�<aAY2+H,���BY1�8t?Ht���at0�2��aA��=�DtvB��O�L_�0��Li�S=��treeview��#X�3��`�381,26�o//A/S/� w/�/�/�/�/�/`/�/ ??+?=?O?�o�
���o%���?�?�?�ADr?>1`��?"2�� GOYOd?v?�_�.E-� �O�O�OxO��@�O0OC_U_g_��6�OF�'_ n_�_�_�_8�_���_ �S�_Qocouo$vo�o 핪o#�oS�o�o 1CUz�os� �����
��y� 3�Z�l�~��������/ ؏���� �2���V� h�z�������?�� ��
��.�@�ϟd�v� ��������M����� �*�<�˯N�r����� ����̿[����&� 8�J�ٿnπϒϤ϶� ��wo�o�ϭo"߉'� E�W�i�{ߎߟ߱��� 1�������/�A�S� e�w�9����������� ��e�>�P�b�t��� ��'��������� ��:L^p��� 5��� $� HZl~��1� ���/ /2/�V/ h/z/�/�/�/?/�/�/ �/
??.?����d?� �?�ߍ�?�?�?�?�? OO)O�?5O_OqO�O �O�O�O�O�O��_&_ 8_J_\_n_�_�/�_�_ �_�_�_�_�_"o4oFo Xojo|oo�o�o�o�o �o�o�o0BTf x������ ��,�>�P�b�t��� ��'���Ώ����� ��:�L�^�p�����C? U?ʟy?�UO�O�#� 5�G�Y�k�~������� ůׯ�����1�C� _z�������¿Կ� �
��.�@�R�d�� �ϚϬϾ�����q�� �*�<�N�`���rߖ� �ߺ���������&� 8�J�\�n��ߒ��� ������{���"�4�F� X�j�|�������������������*de�fault؞*level8a�໯Y�w�! tpst[1]�	��y�tpioG[23���u��d�,>men�u7_l.png�A^13cp5�x]�[4�u6 cp���	//-/?/ ��c/u/�/�/�/�/L/ �/�/??)?;?M?�"�prim=^p�age,74,1�R?�?�?�?�?�?�"�f6class,13�?OO0OBOTO�?�25ZO�O�O�O�O�O�#�<~O_$_6_H_Z_]?o218v?�_�_ �_�_�_�O�26�_o�-o?oQocoB�$U�I_USERVI�EW 1�����R 
���jo䒞o�o=m �o�o	-?�oc u���N��� ���o$�6�H���� ������ˏn���� %�7�I��m������ ��`�ԟ�X�!�3� E�W�i��������ï կx�����/�A�쟿*zoomT�?ZOOMIN�S� 񯺿̿޿�ϥ�&� 8�J�\�n�ϒϤ϶������<*maxr�esn�MAXRES���ω�R�d�v߈� ��=߾��������� *�<�N�`�r�߃�� ���������&�8� ��\�n�������G��� ��������3A ��|����g� �0B�fx ���Y���Q /,/>/P/b//�/�/ �/�/�/q/�/??(? :?�K?Y?k?�/�?�? �?�?�? O�?$O6OHO ZOlOO�O�O�O�O�O �?�O�O	_{OD_V_h_ z_�_/_�_�_�_�_�_ 
o�_.o@oRodovoa